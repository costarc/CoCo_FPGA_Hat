library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
	port(
		cs		: in std_logic;
		A		: in std_logic_vector(15 downto 0);
		D		: out std_logic_vector(7 downto 0)
	);
end rom;

architecture rtl of rom is
type MEMORY is array ( 0 to 8191 ) of std_logic_vector(7 downto 0);
constant rom : MEMORY := (
    x"12",
    x"1a",
    x"50",
    x"10",
    x"ce",
    x"01",
    x"9f",
    x"8e",
    x"00",
    x"00",
    x"6f",
    x"80",
    x"8c",
    x"40",
    x"00",
    x"26",
    x"f9",
    x"86",
    x"7e",
    x"b7",
    x"01",
    x"0c",
    x"8e",
    x"dc",
    x"4d",
    x"bf",
    x"01",
    x"0d",
    x"86",
    x"35",
    x"b7",
    x"ff",
    x"03",
    x"86",
    x"20",
    x"b7",
    x"ff",
    x"98",
    x"86",
    x"fe",
    x"b7",
    x"ff",
    x"02",
    x"b6",
    x"ff",
    x"00",
    x"84",
    x"10",
    x"26",
    x"0f",
    x"cc",
    x"00",
    x"09",
    x"fd",
    x"ff",
    x"b4",
    x"cc",
    x"24",
    x"3f",
    x"fd",
    x"ff",
    x"b6",
    x"86",
    x"e8",
    x"8c",
    x"86",
    x"f8",
    x"97",
    x"6a",
    x"bd",
    x"c2",
    x"01",
    x"cc",
    x"1c",
    x"00",
    x"bd",
    x"cd",
    x"f7",
    x"bd",
    x"cd",
    x"e3",
    x"4f",
    x"bd",
    x"c1",
    x"f6",
    x"bd",
    x"c2",
    x"17",
    x"b7",
    x"ff",
    x"de",
    x"8e",
    x"c0",
    x"00",
    x"9f",
    x"61",
    x"9f",
    x"72",
    x"86",
    x"55",
    x"97",
    x"71",
    x"bd",
    x"db",
    x"ad",
    x"0c",
    x"51",
    x"8e",
    x"03",
    x"6b",
    x"86",
    x"0a",
    x"6f",
    x"80",
    x"4a",
    x"26",
    x"fb",
    x"bd",
    x"dc",
    x"c7",
    x"86",
    x"01",
    x"97",
    x"3a",
    x"bd",
    x"d1",
    x"1a",
    x"86",
    x"0a",
    x"97",
    x"39",
    x"86",
    x"55",
    x"97",
    x"69",
    x"bd",
    x"ce",
    x"0b",
    x"bd",
    x"c2",
    x"01",
    x"cc",
    x"1c",
    x"00",
    x"bd",
    x"cd",
    x"f7",
    x"bd",
    x"cd",
    x"e3",
    x"bd",
    x"ce",
    x"10",
    x"8e",
    x"04",
    x"00",
    x"9f",
    x"4e",
    x"ce",
    x"ce",
    x"c4",
    x"bd",
    x"d2",
    x"4e",
    x"ce",
    x"da",
    x"19",
    x"8e",
    x"c2",
    x"3d",
    x"86",
    x"0d",
    x"97",
    x"26",
    x"34",
    x"10",
    x"ae",
    x"84",
    x"bd",
    x"d8",
    x"e2",
    x"35",
    x"10",
    x"30",
    x"02",
    x"0a",
    x"26",
    x"26",
    x"f1",
    x"ce",
    x"00",
    x"bb",
    x"bd",
    x"c2",
    x"22",
    x"ce",
    x"00",
    x"bb",
    x"8e",
    x"18",
    x"12",
    x"bd",
    x"db",
    x"21",
    x"bd",
    x"d8",
    x"e2",
    x"ce",
    x"00",
    x"c3",
    x"bd",
    x"c2",
    x"22",
    x"ce",
    x"00",
    x"c3",
    x"8e",
    x"19",
    x"52",
    x"bd",
    x"db",
    x"21",
    x"bd",
    x"d8",
    x"e2",
    x"ce",
    x"00",
    x"b3",
    x"8e",
    x"16",
    x"cc",
    x"bd",
    x"db",
    x"21",
    x"bd",
    x"d8",
    x"e2",
    x"cc",
    x"04",
    x"00",
    x"bd",
    x"cd",
    x"f7",
    x"8e",
    x"04",
    x"00",
    x"ec",
    x"84",
    x"ed",
    x"89",
    x"18",
    x"00",
    x"30",
    x"02",
    x"8c",
    x"1c",
    x"00",
    x"26",
    x"f3",
    x"1c",
    x"ef",
    x"96",
    x"51",
    x"97",
    x"50",
    x"86",
    x"01",
    x"97",
    x"52",
    x"bd",
    x"dc",
    x"39",
    x"bd",
    x"dc",
    x"66",
    x"96",
    x"15",
    x"81",
    x"04",
    x"26",
    x"08",
    x"86",
    x"01",
    x"97",
    x"50",
    x"97",
    x"51",
    x"20",
    x"0a",
    x"81",
    x"02",
    x"26",
    x"06",
    x"86",
    x"02",
    x"97",
    x"50",
    x"97",
    x"51",
    x"96",
    x"50",
    x"c6",
    x"ff",
    x"44",
    x"27",
    x"08",
    x"7f",
    x"13",
    x"64",
    x"f7",
    x"13",
    x"70",
    x"20",
    x"06",
    x"f7",
    x"13",
    x"64",
    x"7f",
    x"13",
    x"70",
    x"bd",
    x"cf",
    x"53",
    x"b6",
    x"ff",
    x"00",
    x"85",
    x"01",
    x"26",
    x"c3",
    x"c6",
    x"03",
    x"d7",
    x"55",
    x"d7",
    x"56",
    x"bd",
    x"c2",
    x"0d",
    x"0f",
    x"3a",
    x"86",
    x"01",
    x"97",
    x"52",
    x"ce",
    x"da",
    x"d2",
    x"df",
    x"53",
    x"fc",
    x"d2",
    x"72",
    x"dd",
    x"5e",
    x"0f",
    x"60",
    x"bd",
    x"cb",
    x"a5",
    x"bd",
    x"d1",
    x"1a",
    x"bd",
    x"d1",
    x"4c",
    x"bd",
    x"ce",
    x"b6",
    x"bd",
    x"ce",
    x"cf",
    x"bd",
    x"ce",
    x"fa",
    x"bd",
    x"cc",
    x"a3",
    x"bd",
    x"cc",
    x"d3",
    x"bd",
    x"ce",
    x"68",
    x"10",
    x"8e",
    x"01",
    x"aa",
    x"bd",
    x"c6",
    x"a9",
    x"96",
    x"48",
    x"27",
    x"09",
    x"0f",
    x"48",
    x"10",
    x"8e",
    x"01",
    x"aa",
    x"bd",
    x"d8",
    x"60",
    x"bd",
    x"cc",
    x"b1",
    x"bd",
    x"c3",
    x"b3",
    x"96",
    x"49",
    x"27",
    x"09",
    x"0f",
    x"49",
    x"10",
    x"8e",
    x"01",
    x"bf",
    x"bd",
    x"d8",
    x"60",
    x"8e",
    x"ff",
    x"00",
    x"86",
    x"fb",
    x"a7",
    x"02",
    x"a6",
    x"84",
    x"84",
    x"40",
    x"26",
    x"10",
    x"34",
    x"01",
    x"1a",
    x"50",
    x"86",
    x"fd",
    x"a7",
    x"02",
    x"e6",
    x"84",
    x"c4",
    x"40",
    x"26",
    x"f6",
    x"35",
    x"01",
    x"b6",
    x"01",
    x"a2",
    x"4a",
    x"26",
    x"0e",
    x"b6",
    x"01",
    x"a0",
    x"84",
    x"07",
    x"81",
    x"06",
    x"25",
    x"05",
    x"86",
    x"2f",
    x"b7",
    x"ff",
    x"20",
    x"bd",
    x"cf",
    x"53",
    x"86",
    x"02",
    x"b7",
    x"ff",
    x"20",
    x"bd",
    x"ca",
    x"b6",
    x"bd",
    x"cb",
    x"c3",
    x"96",
    x"14",
    x"27",
    x"04",
    x"0f",
    x"14",
    x"20",
    x"99",
    x"8e",
    x"00",
    x"23",
    x"bd",
    x"dc",
    x"39",
    x"20",
    x"f0",
    x"8e",
    x"7e",
    x"00",
    x"a7",
    x"80",
    x"8c",
    x"80",
    x"00",
    x"26",
    x"f9",
    x"39",
    x"34",
    x"01",
    x"0f",
    x"14",
    x"1c",
    x"ef",
    x"96",
    x"14",
    x"27",
    x"fc",
    x"35",
    x"81",
    x"8e",
    x"00",
    x"bb",
    x"6f",
    x"80",
    x"8c",
    x"00",
    x"d3",
    x"26",
    x"f9",
    x"86",
    x"ff",
    x"97",
    x"ba",
    x"97",
    x"c2",
    x"97",
    x"ca",
    x"97",
    x"d2",
    x"39",
    x"8e",
    x"00",
    x"b3",
    x"34",
    x"50",
    x"a6",
    x"c0",
    x"2b",
    x"06",
    x"a1",
    x"80",
    x"27",
    x"f8",
    x"22",
    x"02",
    x"35",
    x"d0",
    x"35",
    x"50",
    x"a6",
    x"c0",
    x"2b",
    x"e8",
    x"a7",
    x"80",
    x"20",
    x"f8",
    x"07",
    x"c9",
    x"09",
    x"0a",
    x"0a",
    x"47",
    x"0b",
    x"89",
    x"0c",
    x"c6",
    x"0e",
    x"0a",
    x"0f",
    x"47",
    x"10",
    x"86",
    x"13",
    x"05",
    x"13",
    x"11",
    x"15",
    x"8b",
    x"18",
    x"06",
    x"19",
    x"46",
    x"35",
    x"20",
    x"10",
    x"9e",
    x"3d",
    x"86",
    x"0a",
    x"97",
    x"43",
    x"86",
    x"08",
    x"97",
    x"44",
    x"c6",
    x"05",
    x"a6",
    x"a4",
    x"94",
    x"52",
    x"27",
    x"0d",
    x"a6",
    x"22",
    x"dd",
    x"41",
    x"a6",
    x"23",
    x"97",
    x"42",
    x"bd",
    x"c3",
    x"7c",
    x"26",
    x"6b",
    x"31",
    x"25",
    x"5a",
    x"26",
    x"e8",
    x"10",
    x"8e",
    x"01",
    x"ef",
    x"86",
    x"06",
    x"97",
    x"43",
    x"86",
    x"04",
    x"97",
    x"44",
    x"d6",
    x"3f",
    x"a6",
    x"a4",
    x"27",
    x"13",
    x"a6",
    x"23",
    x"97",
    x"41",
    x"a6",
    x"25",
    x"97",
    x"42",
    x"bd",
    x"c3",
    x"7c",
    x"27",
    x"06",
    x"a6",
    x"a4",
    x"2b",
    x"02",
    x"20",
    x"3a",
    x"31",
    x"2d",
    x"5a",
    x"26",
    x"e4",
    x"86",
    x"08",
    x"97",
    x"43",
    x"86",
    x"08",
    x"97",
    x"44",
    x"b6",
    x"01",
    x"c3",
    x"97",
    x"41",
    x"b6",
    x"01",
    x"c5",
    x"97",
    x"42",
    x"bd",
    x"c3",
    x"7c",
    x"26",
    x"1e",
    x"86",
    x"06",
    x"97",
    x"43",
    x"86",
    x"08",
    x"97",
    x"44",
    x"b6",
    x"01",
    x"d8",
    x"97",
    x"41",
    x"b6",
    x"01",
    x"da",
    x"97",
    x"42",
    x"bd",
    x"c3",
    x"7c",
    x"26",
    x"07",
    x"10",
    x"8e",
    x"01",
    x"aa",
    x"7e",
    x"c4",
    x"8c",
    x"10",
    x"8e",
    x"01",
    x"aa",
    x"7e",
    x"c5",
    x"3c",
    x"96",
    x"52",
    x"43",
    x"a4",
    x"a4",
    x"a7",
    x"a4",
    x"e6",
    x"24",
    x"2b",
    x"2c",
    x"8e",
    x"3e",
    x"c0",
    x"30",
    x"85",
    x"a6",
    x"84",
    x"9a",
    x"52",
    x"a7",
    x"84",
    x"bd",
    x"cc",
    x"a7",
    x"e1",
    x"05",
    x"27",
    x"0a",
    x"30",
    x"89",
    x"00",
    x"06",
    x"a6",
    x"84",
    x"26",
    x"f4",
    x"20",
    x"10",
    x"ce",
    x"1c",
    x"00",
    x"df",
    x"4e",
    x"bd",
    x"cd",
    x"81",
    x"ce",
    x"04",
    x"00",
    x"df",
    x"4e",
    x"bd",
    x"cd",
    x"81",
    x"dc",
    x"1b",
    x"bd",
    x"dc",
    x"39",
    x"c4",
    x"7f",
    x"a6",
    x"21",
    x"27",
    x"0e",
    x"4a",
    x"27",
    x"06",
    x"4f",
    x"c3",
    x"00",
    x"c8",
    x"20",
    x"08",
    x"c3",
    x"01",
    x"2c",
    x"20",
    x"03",
    x"c3",
    x"01",
    x"90",
    x"34",
    x"20",
    x"bd",
    x"db",
    x"0c",
    x"35",
    x"20",
    x"bd",
    x"d1",
    x"42",
    x"d7",
    x"26",
    x"8d",
    x"0c",
    x"cc",
    x"12",
    x"80",
    x"8d",
    x"15",
    x"10",
    x"8e",
    x"01",
    x"aa",
    x"7e",
    x"d8",
    x"60",
    x"ec",
    x"89",
    x"18",
    x"00",
    x"ed",
    x"84",
    x"30",
    x"88",
    x"20",
    x"0a",
    x"26",
    x"26",
    x"f3",
    x"39",
    x"97",
    x"4d",
    x"d7",
    x"26",
    x"86",
    x"ff",
    x"b7",
    x"ff",
    x"20",
    x"8d",
    x"0c",
    x"86",
    x"02",
    x"b7",
    x"ff",
    x"20",
    x"8d",
    x"05",
    x"0a",
    x"26",
    x"26",
    x"ee",
    x"39",
    x"d6",
    x"4d",
    x"5a",
    x"26",
    x"fd",
    x"39",
    x"8e",
    x"01",
    x"aa",
    x"a6",
    x"04",
    x"91",
    x"41",
    x"23",
    x"08",
    x"90",
    x"41",
    x"91",
    x"43",
    x"23",
    x"0a",
    x"20",
    x"20",
    x"96",
    x"41",
    x"a0",
    x"04",
    x"a1",
    x"1f",
    x"22",
    x"18",
    x"a6",
    x"06",
    x"91",
    x"42",
    x"23",
    x"08",
    x"90",
    x"42",
    x"91",
    x"44",
    x"23",
    x"0e",
    x"20",
    x"0a",
    x"96",
    x"42",
    x"a0",
    x"06",
    x"81",
    x"08",
    x"23",
    x"04",
    x"20",
    x"00",
    x"4f",
    x"39",
    x"86",
    x"ff",
    x"39",
    x"39",
    x"10",
    x"8e",
    x"01",
    x"aa",
    x"a6",
    x"38",
    x"4a",
    x"26",
    x"05",
    x"c6",
    x"3f",
    x"f7",
    x"ff",
    x"20",
    x"a6",
    x"3b",
    x"27",
    x"ed",
    x"81",
    x"01",
    x"10",
    x"27",
    x"00",
    x"c1",
    x"96",
    x"30",
    x"10",
    x"26",
    x"01",
    x"7b",
    x"a6",
    x"3e",
    x"10",
    x"2b",
    x"02",
    x"e1",
    x"10",
    x"26",
    x"00",
    x"bd",
    x"6c",
    x"36",
    x"ce",
    x"3b",
    x"80",
    x"a6",
    x"38",
    x"c6",
    x"3c",
    x"3d",
    x"33",
    x"cb",
    x"a6",
    x"26",
    x"84",
    x"03",
    x"c6",
    x"0f",
    x"3d",
    x"33",
    x"cb",
    x"a6",
    x"38",
    x"81",
    x"03",
    x"22",
    x"08",
    x"a6",
    x"3c",
    x"26",
    x"04",
    x"33",
    x"c9",
    x"01",
    x"68",
    x"ae",
    x"2c",
    x"30",
    x"88",
    x"20",
    x"34",
    x"20",
    x"10",
    x"8e",
    x"00",
    x"74",
    x"86",
    x"05",
    x"97",
    x"26",
    x"37",
    x"06",
    x"a4",
    x"84",
    x"aa",
    x"89",
    x"18",
    x"00",
    x"a7",
    x"a0",
    x"e4",
    x"01",
    x"ea",
    x"89",
    x"18",
    x"01",
    x"e7",
    x"a0",
    x"37",
    x"02",
    x"a4",
    x"02",
    x"aa",
    x"89",
    x"18",
    x"02",
    x"a7",
    x"a0",
    x"30",
    x"88",
    x"60",
    x"0a",
    x"26",
    x"26",
    x"dd",
    x"35",
    x"20",
    x"ce",
    x"34",
    x"00",
    x"a6",
    x"38",
    x"c6",
    x"c0",
    x"3d",
    x"33",
    x"cb",
    x"a6",
    x"26",
    x"84",
    x"03",
    x"c6",
    x"30",
    x"3d",
    x"33",
    x"cb",
    x"33",
    x"43",
    x"a6",
    x"38",
    x"81",
    x"03",
    x"22",
    x"08",
    x"a6",
    x"3c",
    x"26",
    x"04",
    x"33",
    x"c9",
    x"04",
    x"80",
    x"ae",
    x"2c",
    x"30",
    x"89",
    x"18",
    x"20",
    x"34",
    x"20",
    x"10",
    x"8e",
    x"00",
    x"74",
    x"86",
    x"05",
    x"97",
    x"26",
    x"37",
    x"06",
    x"aa",
    x"84",
    x"a1",
    x"a0",
    x"10",
    x"26",
    x"fd",
    x"e8",
    x"ea",
    x"01",
    x"e1",
    x"a0",
    x"10",
    x"26",
    x"fd",
    x"e0",
    x"37",
    x"02",
    x"aa",
    x"02",
    x"a1",
    x"a0",
    x"10",
    x"26",
    x"fd",
    x"d6",
    x"30",
    x"88",
    x"60",
    x"33",
    x"46",
    x"0a",
    x"26",
    x"26",
    x"db",
    x"35",
    x"20",
    x"96",
    x"2c",
    x"10",
    x"26",
    x"03",
    x"17",
    x"a6",
    x"35",
    x"10",
    x"26",
    x"00",
    x"94",
    x"8d",
    x"4d",
    x"30",
    x"89",
    x"02",
    x"00",
    x"ce",
    x"c5",
    x"0d",
    x"ec",
    x"c6",
    x"a4",
    x"89",
    x"18",
    x"00",
    x"e4",
    x"89",
    x"18",
    x"01",
    x"10",
    x"93",
    x"1b",
    x"27",
    x"0e",
    x"34",
    x"04",
    x"bd",
    x"ca",
    x"9b",
    x"35",
    x"02",
    x"26",
    x"73",
    x"bd",
    x"ca",
    x"9b",
    x"26",
    x"6e",
    x"86",
    x"ff",
    x"97",
    x"2d",
    x"ec",
    x"a4",
    x"c3",
    x"00",
    x"06",
    x"10",
    x"83",
    x"01",
    x"00",
    x"23",
    x"05",
    x"0f",
    x"2e",
    x"cc",
    x"01",
    x"00",
    x"ed",
    x"a4",
    x"96",
    x"2e",
    x"2b",
    x"2a",
    x"a6",
    x"3c",
    x"2b",
    x"1b",
    x"ec",
    x"22",
    x"c3",
    x"00",
    x"01",
    x"2b",
    x"1d",
    x"dc",
    x"1b",
    x"20",
    x"19",
    x"8e",
    x"c5",
    x"09",
    x"e6",
    x"26",
    x"c4",
    x"03",
    x"1f",
    x"98",
    x"e6",
    x"85",
    x"ae",
    x"28",
    x"3a",
    x"48",
    x"39",
    x"ec",
    x"22",
    x"c3",
    x"ff",
    x"ff",
    x"2a",
    x"02",
    x"dc",
    x"1b",
    x"ed",
    x"22",
    x"a6",
    x"3e",
    x"26",
    x"69",
    x"7e",
    x"c7",
    x"83",
    x"00",
    x"00",
    x"00",
    x"01",
    x"03",
    x"c0",
    x"00",
    x"f0",
    x"00",
    x"3c",
    x"0f",
    x"00",
    x"3f",
    x"f0",
    x"0f",
    x"fc",
    x"03",
    x"ff",
    x"ff",
    x"c0",
    x"03",
    x"00",
    x"00",
    x"c0",
    x"00",
    x"30",
    x"0c",
    x"00",
    x"dc",
    x"1b",
    x"ed",
    x"a4",
    x"ed",
    x"22",
    x"39",
    x"0f",
    x"2d",
    x"a6",
    x"3e",
    x"26",
    x"3d",
    x"ec",
    x"a4",
    x"10",
    x"83",
    x"01",
    x"00",
    x"10",
    x"26",
    x"01",
    x"dc",
    x"8d",
    x"e7",
    x"6f",
    x"35",
    x"0f",
    x"2c",
    x"0f",
    x"2f",
    x"96",
    x"2d",
    x"27",
    x"1c",
    x"86",
    x"32",
    x"97",
    x"30",
    x"0a",
    x"30",
    x"27",
    x"14",
    x"96",
    x"30",
    x"84",
    x"04",
    x"27",
    x"05",
    x"86",
    x"ff",
    x"a7",
    x"3c",
    x"8c",
    x"6f",
    x"3c",
    x"86",
    x"02",
    x"a7",
    x"38",
    x"7e",
    x"c9",
    x"7f",
    x"86",
    x"0a",
    x"a7",
    x"3d",
    x"86",
    x"02",
    x"a7",
    x"3e",
    x"7e",
    x"c3",
    x"b2",
    x"96",
    x"2d",
    x"26",
    x"93",
    x"8d",
    x"b0",
    x"a6",
    x"3e",
    x"4a",
    x"27",
    x"32",
    x"8e",
    x"00",
    x"83",
    x"86",
    x"30",
    x"6f",
    x"80",
    x"4a",
    x"26",
    x"fb",
    x"8e",
    x"00",
    x"98",
    x"ce",
    x"de",
    x"ef",
    x"86",
    x"1b",
    x"e6",
    x"c0",
    x"e7",
    x"80",
    x"4a",
    x"26",
    x"f9",
    x"a6",
    x"26",
    x"84",
    x"03",
    x"27",
    x"07",
    x"97",
    x"26",
    x"c6",
    x"10",
    x"bd",
    x"cd",
    x"c9",
    x"cc",
    x"25",
    x"08",
    x"bd",
    x"c3",
    x"5f",
    x"ce",
    x"00",
    x"83",
    x"bd",
    x"c9",
    x"a2",
    x"6a",
    x"3d",
    x"10",
    x"26",
    x"fe",
    x"00",
    x"6a",
    x"3e",
    x"27",
    x"28",
    x"86",
    x"0c",
    x"a7",
    x"3f",
    x"17",
    x"12",
    x"f8",
    x"86",
    x"10",
    x"a7",
    x"3f",
    x"86",
    x"46",
    x"a7",
    x"3d",
    x"16",
    x"fd",
    x"ea",
    x"8e",
    x"c5",
    x"d2",
    x"96",
    x"52",
    x"84",
    x"02",
    x"ae",
    x"86",
    x"39",
    x"00",
    x"55",
    x"00",
    x"56",
    x"00",
    x"57",
    x"00",
    x"5c",
    x"da",
    x"da",
    x"da",
    x"ef",
    x"b6",
    x"01",
    x"cf",
    x"27",
    x"11",
    x"bd",
    x"cb",
    x"b9",
    x"d6",
    x"39",
    x"58",
    x"3a",
    x"cc",
    x"08",
    x"00",
    x"ed",
    x"84",
    x"86",
    x"ff",
    x"b7",
    x"01",
    x"cf",
    x"8d",
    x"d2",
    x"a6",
    x"84",
    x"81",
    x"05",
    x"23",
    x"04",
    x"86",
    x"05",
    x"a7",
    x"84",
    x"6a",
    x"84",
    x"10",
    x"2b",
    x"16",
    x"06",
    x"34",
    x"20",
    x"96",
    x"50",
    x"84",
    x"02",
    x"10",
    x"27",
    x"00",
    x"95",
    x"96",
    x"52",
    x"84",
    x"02",
    x"26",
    x"0a",
    x"0c",
    x"52",
    x"ce",
    x"da",
    x"d6",
    x"8e",
    x"00",
    x"57",
    x"20",
    x"08",
    x"0a",
    x"52",
    x"ce",
    x"da",
    x"d2",
    x"8e",
    x"00",
    x"5c",
    x"df",
    x"53",
    x"a6",
    x"24",
    x"e6",
    x"26",
    x"ed",
    x"02",
    x"96",
    x"39",
    x"a7",
    x"04",
    x"bd",
    x"ce",
    x"10",
    x"cc",
    x"1c",
    x"00",
    x"bd",
    x"cd",
    x"f7",
    x"ce",
    x"ce",
    x"c4",
    x"bd",
    x"d2",
    x"4e",
    x"96",
    x"52",
    x"84",
    x"02",
    x"8e",
    x"c5",
    x"da",
    x"ee",
    x"86",
    x"8e",
    x"0f",
    x"66",
    x"bd",
    x"d8",
    x"e2",
    x"bd",
    x"c2",
    x"01",
    x"1c",
    x"ef",
    x"cc",
    x"04",
    x"00",
    x"bd",
    x"cd",
    x"f7",
    x"8e",
    x"04",
    x"00",
    x"ec",
    x"81",
    x"ed",
    x"89",
    x"17",
    x"fe",
    x"8c",
    x"1c",
    x"00",
    x"26",
    x"f5",
    x"bd",
    x"d1",
    x"1a",
    x"86",
    x"0a",
    x"97",
    x"3f",
    x"97",
    x"39",
    x"bd",
    x"cf",
    x"53",
    x"8e",
    x"ff",
    x"00",
    x"86",
    x"ff",
    x"a7",
    x"02",
    x"a6",
    x"84",
    x"95",
    x"52",
    x"27",
    x"12",
    x"85",
    x"01",
    x"27",
    x"ec",
    x"85",
    x"02",
    x"27",
    x"e8",
    x"6f",
    x"02",
    x"a6",
    x"84",
    x"8a",
    x"83",
    x"81",
    x"ff",
    x"27",
    x"de",
    x"8e",
    x"c5",
    x"d6",
    x"96",
    x"52",
    x"84",
    x"02",
    x"ae",
    x"86",
    x"10",
    x"ae",
    x"e4",
    x"bd",
    x"cc",
    x"d3",
    x"35",
    x"20",
    x"6c",
    x"3b",
    x"86",
    x"28",
    x"a7",
    x"3d",
    x"cc",
    x"01",
    x"90",
    x"dd",
    x"4b",
    x"86",
    x"ff",
    x"a7",
    x"3e",
    x"6f",
    x"38",
    x"bd",
    x"dc",
    x"66",
    x"96",
    x"15",
    x"27",
    x"04",
    x"dc",
    x"1b",
    x"dd",
    x"4b",
    x"4f",
    x"dc",
    x"4b",
    x"27",
    x"05",
    x"83",
    x"00",
    x"01",
    x"dd",
    x"4b",
    x"a6",
    x"3d",
    x"27",
    x"03",
    x"4a",
    x"a7",
    x"3d",
    x"26",
    x"5a",
    x"dc",
    x"4b",
    x"26",
    x"56",
    x"34",
    x"20",
    x"10",
    x"8e",
    x"01",
    x"e9",
    x"bd",
    x"c5",
    x"c8",
    x"a6",
    x"84",
    x"e6",
    x"3b",
    x"3d",
    x"ae",
    x"22",
    x"30",
    x"8b",
    x"a6",
    x"3f",
    x"97",
    x"26",
    x"dc",
    x"1b",
    x"ed",
    x"84",
    x"30",
    x"88",
    x"20",
    x"0a",
    x"26",
    x"26",
    x"f7",
    x"35",
    x"20",
    x"6f",
    x"3e",
    x"ae",
    x"28",
    x"e6",
    x"3f",
    x"d7",
    x"26",
    x"ec",
    x"89",
    x"18",
    x"00",
    x"ed",
    x"84",
    x"a6",
    x"89",
    x"18",
    x"02",
    x"a7",
    x"02",
    x"30",
    x"88",
    x"20",
    x"0a",
    x"26",
    x"26",
    x"ed",
    x"a6",
    x"35",
    x"2b",
    x"18",
    x"ec",
    x"a4",
    x"27",
    x"14",
    x"86",
    x"04",
    x"97",
    x"2f",
    x"6f",
    x"38",
    x"0f",
    x"2e",
    x"86",
    x"7f",
    x"b7",
    x"ff",
    x"20",
    x"7e",
    x"c7",
    x"be",
    x"4f",
    x"7e",
    x"c8",
    x"5f",
    x"bd",
    x"dc",
    x"66",
    x"a6",
    x"35",
    x"27",
    x"28",
    x"81",
    x"01",
    x"10",
    x"27",
    x"00",
    x"86",
    x"96",
    x"15",
    x"81",
    x"02",
    x"27",
    x"13",
    x"81",
    x"04",
    x"27",
    x"08",
    x"0f",
    x"2c",
    x"0f",
    x"2f",
    x"0f",
    x"2e",
    x"20",
    x"74",
    x"6f",
    x"3c",
    x"cc",
    x"ff",
    x"ca",
    x"20",
    x"07",
    x"86",
    x"ff",
    x"a7",
    x"3c",
    x"cc",
    x"00",
    x"36",
    x"ed",
    x"22",
    x"96",
    x"52",
    x"b5",
    x"ff",
    x"00",
    x"26",
    x"5d",
    x"96",
    x"31",
    x"26",
    x"5b",
    x"0a",
    x"31",
    x"96",
    x"2f",
    x"26",
    x"53",
    x"cc",
    x"ff",
    x"61",
    x"ed",
    x"a4",
    x"86",
    x"28",
    x"97",
    x"2c",
    x"86",
    x"ff",
    x"97",
    x"2e",
    x"97",
    x"2d",
    x"7e",
    x"c8",
    x"6f",
    x"e6",
    x"26",
    x"a6",
    x"3c",
    x"27",
    x"04",
    x"cb",
    x"04",
    x"20",
    x"02",
    x"c0",
    x"04",
    x"e7",
    x"26",
    x"bd",
    x"c5",
    x"25",
    x"97",
    x"36",
    x"a6",
    x"35",
    x"2b",
    x"05",
    x"6f",
    x"35",
    x"7e",
    x"c8",
    x"79",
    x"86",
    x"01",
    x"a7",
    x"35",
    x"7e",
    x"c8",
    x"79",
    x"96",
    x"2c",
    x"48",
    x"8a",
    x"02",
    x"b7",
    x"ff",
    x"20",
    x"ec",
    x"a4",
    x"c3",
    x"00",
    x"03",
    x"ed",
    x"a4",
    x"0a",
    x"2c",
    x"10",
    x"26",
    x"00",
    x"bb",
    x"dc",
    x"1b",
    x"ed",
    x"a4",
    x"a7",
    x"35",
    x"7e",
    x"c8",
    x"79",
    x"0f",
    x"31",
    x"96",
    x"15",
    x"10",
    x"2b",
    x"00",
    x"8a",
    x"27",
    x"39",
    x"81",
    x"02",
    x"25",
    x"28",
    x"27",
    x"5e",
    x"81",
    x"03",
    x"27",
    x"42",
    x"a6",
    x"3c",
    x"27",
    x"04",
    x"0f",
    x"36",
    x"6f",
    x"3c",
    x"a6",
    x"35",
    x"27",
    x"0f",
    x"bd",
    x"c5",
    x"25",
    x"0c",
    x"36",
    x"96",
    x"36",
    x"81",
    x"14",
    x"22",
    x"94",
    x"dc",
    x"1b",
    x"20",
    x"03",
    x"cc",
    x"ff",
    x"ca",
    x"ed",
    x"22",
    x"20",
    x"5c",
    x"0f",
    x"36",
    x"a6",
    x"35",
    x"2a",
    x"07",
    x"cc",
    x"ff",
    x"c0",
    x"ed",
    x"a4",
    x"20",
    x"1e",
    x"0f",
    x"36",
    x"bd",
    x"c5",
    x"25",
    x"e6",
    x"35",
    x"2a",
    x"4c",
    x"a6",
    x"38",
    x"81",
    x"03",
    x"22",
    x"02",
    x"86",
    x"04",
    x"20",
    x"14",
    x"0f",
    x"36",
    x"a6",
    x"35",
    x"2a",
    x"e7",
    x"cc",
    x"00",
    x"70",
    x"ed",
    x"a4",
    x"a6",
    x"36",
    x"44",
    x"44",
    x"44",
    x"84",
    x"01",
    x"8b",
    x"04",
    x"a7",
    x"38",
    x"20",
    x"44",
    x"a6",
    x"3c",
    x"2b",
    x"06",
    x"0f",
    x"36",
    x"86",
    x"ff",
    x"a7",
    x"3c",
    x"a6",
    x"35",
    x"27",
    x"11",
    x"bd",
    x"c5",
    x"25",
    x"0c",
    x"36",
    x"96",
    x"36",
    x"81",
    x"14",
    x"10",
    x"22",
    x"ff",
    x"36",
    x"dc",
    x"1b",
    x"20",
    x"03",
    x"cc",
    x"00",
    x"36",
    x"ed",
    x"22",
    x"a6",
    x"36",
    x"44",
    x"44",
    x"84",
    x"03",
    x"e6",
    x"35",
    x"27",
    x"0e",
    x"2a",
    x"0a",
    x"a6",
    x"38",
    x"81",
    x"03",
    x"22",
    x"06",
    x"86",
    x"05",
    x"20",
    x"02",
    x"86",
    x"02",
    x"a7",
    x"38",
    x"d6",
    x"2f",
    x"27",
    x"02",
    x"0a",
    x"2f",
    x"a6",
    x"35",
    x"81",
    x"01",
    x"27",
    x"78",
    x"bd",
    x"c4",
    x"e7",
    x"30",
    x"89",
    x"01",
    x"00",
    x"ce",
    x"c5",
    x"1d",
    x"ec",
    x"c6",
    x"a4",
    x"89",
    x"18",
    x"00",
    x"e4",
    x"89",
    x"18",
    x"01",
    x"10",
    x"93",
    x"1b",
    x"27",
    x"1d",
    x"34",
    x"04",
    x"8d",
    x"1d",
    x"35",
    x"02",
    x"26",
    x"04",
    x"8d",
    x"17",
    x"27",
    x"11",
    x"a6",
    x"35",
    x"2b",
    x"1a",
    x"86",
    x"ff",
    x"a7",
    x"35",
    x"bd",
    x"c5",
    x"25",
    x"0f",
    x"2c",
    x"0f",
    x"2e",
    x"20",
    x"0d",
    x"6f",
    x"35",
    x"20",
    x"3e",
    x"bd",
    x"ca",
    x"9b",
    x"96",
    x"4d",
    x"43",
    x"94",
    x"34",
    x"39",
    x"96",
    x"2c",
    x"26",
    x"31",
    x"ec",
    x"a4",
    x"2a",
    x"2d",
    x"bd",
    x"c4",
    x"e7",
    x"30",
    x"89",
    x"00",
    x"e0",
    x"ce",
    x"c5",
    x"1d",
    x"ec",
    x"c6",
    x"a4",
    x"89",
    x"18",
    x"00",
    x"e4",
    x"89",
    x"18",
    x"01",
    x"10",
    x"93",
    x"1b",
    x"27",
    x"0c",
    x"34",
    x"04",
    x"8d",
    x"d2",
    x"35",
    x"02",
    x"26",
    x"0c",
    x"8d",
    x"cc",
    x"26",
    x"08",
    x"86",
    x"04",
    x"a7",
    x"38",
    x"dc",
    x"1b",
    x"ed",
    x"a4",
    x"ec",
    x"24",
    x"e3",
    x"a4",
    x"ed",
    x"24",
    x"ec",
    x"26",
    x"e3",
    x"22",
    x"ed",
    x"26",
    x"a6",
    x"35",
    x"27",
    x"12",
    x"96",
    x"23",
    x"a1",
    x"24",
    x"27",
    x"0c",
    x"a6",
    x"36",
    x"84",
    x"07",
    x"48",
    x"48",
    x"48",
    x"8a",
    x"1a",
    x"b7",
    x"ff",
    x"20",
    x"a6",
    x"24",
    x"97",
    x"23",
    x"a6",
    x"35",
    x"26",
    x"59",
    x"8e",
    x"c5",
    x"09",
    x"e6",
    x"26",
    x"c4",
    x"03",
    x"1f",
    x"98",
    x"e6",
    x"85",
    x"34",
    x"06",
    x"bd",
    x"d8",
    x"52",
    x"ed",
    x"28",
    x"1f",
    x"01",
    x"35",
    x"06",
    x"30",
    x"89",
    x"01",
    x"e0",
    x"3a",
    x"48",
    x"ce",
    x"c5",
    x"0d",
    x"ec",
    x"c6",
    x"a4",
    x"89",
    x"18",
    x"00",
    x"e4",
    x"89",
    x"18",
    x"01",
    x"10",
    x"93",
    x"1b",
    x"27",
    x"30",
    x"34",
    x"04",
    x"bd",
    x"ca",
    x"9b",
    x"35",
    x"02",
    x"26",
    x"05",
    x"bd",
    x"ca",
    x"9b",
    x"27",
    x"22",
    x"ec",
    x"26",
    x"a3",
    x"22",
    x"ed",
    x"26",
    x"96",
    x"2c",
    x"26",
    x"04",
    x"6f",
    x"38",
    x"20",
    x"0f",
    x"86",
    x"01",
    x"97",
    x"2c",
    x"ec",
    x"22",
    x"43",
    x"53",
    x"c3",
    x"00",
    x"01",
    x"ed",
    x"22",
    x"63",
    x"3c",
    x"bd",
    x"d8",
    x"52",
    x"ed",
    x"28",
    x"ce",
    x"34",
    x"00",
    x"a6",
    x"38",
    x"81",
    x"03",
    x"22",
    x"08",
    x"a6",
    x"3c",
    x"26",
    x"04",
    x"33",
    x"c9",
    x"04",
    x"80",
    x"a6",
    x"38",
    x"c6",
    x"c0",
    x"3d",
    x"33",
    x"cb",
    x"df",
    x"37",
    x"a6",
    x"26",
    x"84",
    x"03",
    x"c6",
    x"30",
    x"3d",
    x"33",
    x"cb",
    x"ef",
    x"2a",
    x"11",
    x"a3",
    x"2e",
    x"26",
    x"10",
    x"a6",
    x"3e",
    x"2b",
    x"0c",
    x"ee",
    x"28",
    x"11",
    x"a3",
    x"2c",
    x"10",
    x"27",
    x"f9",
    x"fc",
    x"0c",
    x"48",
    x"39",
    x"a6",
    x"3e",
    x"10",
    x"2e",
    x"00",
    x"d9",
    x"e6",
    x"3c",
    x"34",
    x"20",
    x"10",
    x"8e",
    x"01",
    x"e9",
    x"a7",
    x"3e",
    x"e7",
    x"3c",
    x"de",
    x"37",
    x"ef",
    x"a4",
    x"ee",
    x"22",
    x"ef",
    x"24",
    x"bd",
    x"c5",
    x"c8",
    x"a6",
    x"84",
    x"e6",
    x"3e",
    x"2a",
    x"01",
    x"4c",
    x"a7",
    x"3d",
    x"20",
    x"02",
    x"6a",
    x"3d",
    x"10",
    x"27",
    x"00",
    x"af",
    x"ae",
    x"24",
    x"ee",
    x"a4",
    x"a6",
    x"3f",
    x"97",
    x"26",
    x"a6",
    x"3e",
    x"10",
    x"2a",
    x"00",
    x"87",
    x"a6",
    x"3d",
    x"81",
    x"01",
    x"10",
    x"26",
    x"00",
    x"7f",
    x"ce",
    x"34",
    x"00",
    x"a6",
    x"3c",
    x"26",
    x"04",
    x"33",
    x"c9",
    x"04",
    x"80",
    x"df",
    x"45",
    x"bd",
    x"dc",
    x"39",
    x"1f",
    x"52",
    x"31",
    x"a5",
    x"ec",
    x"c4",
    x"48",
    x"58",
    x"aa",
    x"c0",
    x"ea",
    x"c0",
    x"a4",
    x"a0",
    x"e4",
    x"a0",
    x"ed",
    x"84",
    x"a6",
    x"c4",
    x"48",
    x"aa",
    x"c0",
    x"a4",
    x"a0",
    x"a7",
    x"02",
    x"30",
    x"88",
    x"20",
    x"0a",
    x"26",
    x"26",
    x"e2",
    x"10",
    x"8e",
    x"01",
    x"aa",
    x"ae",
    x"28",
    x"af",
    x"2c",
    x"a6",
    x"3f",
    x"97",
    x"26",
    x"de",
    x"45",
    x"a6",
    x"26",
    x"84",
    x"03",
    x"c6",
    x"30",
    x"3d",
    x"33",
    x"cb",
    x"6f",
    x"2e",
    x"bd",
    x"dc",
    x"39",
    x"1f",
    x"52",
    x"31",
    x"a5",
    x"ec",
    x"c4",
    x"48",
    x"58",
    x"aa",
    x"c0",
    x"ea",
    x"c0",
    x"a4",
    x"a0",
    x"aa",
    x"89",
    x"18",
    x"00",
    x"e4",
    x"a0",
    x"ea",
    x"89",
    x"18",
    x"01",
    x"ed",
    x"84",
    x"a6",
    x"c4",
    x"48",
    x"aa",
    x"c0",
    x"a4",
    x"a0",
    x"aa",
    x"89",
    x"18",
    x"02",
    x"a7",
    x"02",
    x"30",
    x"88",
    x"20",
    x"0a",
    x"26",
    x"26",
    x"d6",
    x"35",
    x"20",
    x"39",
    x"37",
    x"06",
    x"ed",
    x"84",
    x"37",
    x"02",
    x"a7",
    x"02",
    x"30",
    x"88",
    x"20",
    x"0a",
    x"26",
    x"26",
    x"f1",
    x"ae",
    x"24",
    x"a6",
    x"3b",
    x"30",
    x"86",
    x"af",
    x"24",
    x"7e",
    x"c9",
    x"e1",
    x"35",
    x"20",
    x"0c",
    x"48",
    x"39",
    x"97",
    x"34",
    x"84",
    x"55",
    x"48",
    x"97",
    x"35",
    x"96",
    x"34",
    x"84",
    x"aa",
    x"44",
    x"9a",
    x"35",
    x"98",
    x"34",
    x"97",
    x"4d",
    x"94",
    x"34",
    x"84",
    x"55",
    x"39",
    x"7e",
    x"ce",
    x"75",
    x"39",
    x"10",
    x"8e",
    x"01",
    x"bf",
    x"a6",
    x"3b",
    x"27",
    x"f4",
    x"96",
    x"32",
    x"2e",
    x"70",
    x"2b",
    x"5f",
    x"8e",
    x"c5",
    x"09",
    x"e6",
    x"26",
    x"c4",
    x"03",
    x"1f",
    x"98",
    x"e6",
    x"85",
    x"ae",
    x"28",
    x"30",
    x"89",
    x"01",
    x"00",
    x"3a",
    x"48",
    x"ce",
    x"cb",
    x"10",
    x"ec",
    x"c6",
    x"a4",
    x"89",
    x"18",
    x"00",
    x"e4",
    x"89",
    x"18",
    x"01",
    x"10",
    x"93",
    x"1b",
    x"27",
    x"0c",
    x"34",
    x"04",
    x"8d",
    x"ae",
    x"35",
    x"02",
    x"26",
    x"27",
    x"8d",
    x"a8",
    x"26",
    x"23",
    x"ec",
    x"a4",
    x"c3",
    x"00",
    x"12",
    x"10",
    x"83",
    x"01",
    x"00",
    x"23",
    x"03",
    x"cc",
    x"01",
    x"00",
    x"ed",
    x"a4",
    x"a6",
    x"3e",
    x"81",
    x"0a",
    x"24",
    x"03",
    x"4c",
    x"a7",
    x"3e",
    x"20",
    x"31",
    x"03",
    x"00",
    x"00",
    x"c0",
    x"00",
    x"30",
    x"0c",
    x"00",
    x"cc",
    x"ff",
    x"00",
    x"ed",
    x"a4",
    x"86",
    x"fb",
    x"97",
    x"32",
    x"20",
    x"6a",
    x"0c",
    x"32",
    x"2b",
    x"66",
    x"cc",
    x"ff",
    x"00",
    x"ed",
    x"a4",
    x"86",
    x"0a",
    x"97",
    x"32",
    x"20",
    x"0f",
    x"ec",
    x"a4",
    x"c3",
    x"00",
    x"0a",
    x"ed",
    x"a4",
    x"0a",
    x"32",
    x"26",
    x"04",
    x"dc",
    x"1b",
    x"ed",
    x"a4",
    x"ec",
    x"24",
    x"e3",
    x"a4",
    x"ed",
    x"24",
    x"ec",
    x"26",
    x"e3",
    x"22",
    x"ed",
    x"26",
    x"8e",
    x"c5",
    x"09",
    x"e6",
    x"26",
    x"c4",
    x"03",
    x"1f",
    x"98",
    x"e6",
    x"85",
    x"34",
    x"06",
    x"bd",
    x"d8",
    x"52",
    x"ed",
    x"28",
    x"1f",
    x"01",
    x"35",
    x"06",
    x"30",
    x"89",
    x"00",
    x"a0",
    x"3a",
    x"48",
    x"ce",
    x"c5",
    x"15",
    x"ec",
    x"c6",
    x"a4",
    x"89",
    x"18",
    x"00",
    x"e4",
    x"89",
    x"18",
    x"01",
    x"10",
    x"93",
    x"1b",
    x"27",
    x"12",
    x"34",
    x"04",
    x"bd",
    x"ca",
    x"9b",
    x"35",
    x"02",
    x"26",
    x"05",
    x"bd",
    x"ca",
    x"9b",
    x"27",
    x"04",
    x"86",
    x"ff",
    x"a7",
    x"3b",
    x"ce",
    x"3d",
    x"d8",
    x"96",
    x"32",
    x"2a",
    x"03",
    x"33",
    x"c8",
    x"60",
    x"a6",
    x"26",
    x"84",
    x"03",
    x"c6",
    x"18",
    x"3d",
    x"33",
    x"cb",
    x"ef",
    x"2a",
    x"0c",
    x"49",
    x"39",
    x"8d",
    x"12",
    x"c6",
    x"14",
    x"d7",
    x"26",
    x"cc",
    x"10",
    x"00",
    x"ed",
    x"81",
    x"0a",
    x"26",
    x"26",
    x"fa",
    x"39",
    x"3e",
    x"98",
    x"3e",
    x"ac",
    x"8e",
    x"cb",
    x"b5",
    x"96",
    x"52",
    x"84",
    x"02",
    x"ae",
    x"86",
    x"39",
    x"d6",
    x"39",
    x"58",
    x"8d",
    x"f1",
    x"ec",
    x"85",
    x"8e",
    x"1b",
    x"14",
    x"bd",
    x"db",
    x"36",
    x"8d",
    x"e7",
    x"0f",
    x"26",
    x"d6",
    x"26",
    x"c1",
    x"0a",
    x"27",
    x"1a",
    x"d1",
    x"39",
    x"27",
    x"10",
    x"ec",
    x"84",
    x"c3",
    x"00",
    x"01",
    x"10",
    x"83",
    x"10",
    x"00",
    x"23",
    x"03",
    x"cc",
    x"10",
    x"00",
    x"ed",
    x"84",
    x"30",
    x"02",
    x"0c",
    x"26",
    x"20",
    x"e0",
    x"10",
    x"8e",
    x"01",
    x"d4",
    x"a6",
    x"3b",
    x"26",
    x"39",
    x"b6",
    x"01",
    x"a8",
    x"2b",
    x"11",
    x"8d",
    x"b6",
    x"d6",
    x"39",
    x"58",
    x"3a",
    x"ec",
    x"84",
    x"27",
    x"0a",
    x"83",
    x"00",
    x"01",
    x"27",
    x"03",
    x"ed",
    x"84",
    x"39",
    x"ed",
    x"84",
    x"cc",
    x"1a",
    x"23",
    x"a7",
    x"24",
    x"e7",
    x"26",
    x"bd",
    x"d8",
    x"52",
    x"ed",
    x"28",
    x"86",
    x"01",
    x"a7",
    x"3b",
    x"86",
    x"06",
    x"a7",
    x"3f",
    x"86",
    x"01",
    x"bd",
    x"dc",
    x"39",
    x"ed",
    x"a4",
    x"bd",
    x"dc",
    x"39",
    x"ed",
    x"22",
    x"6c",
    x"3d",
    x"a6",
    x"3d",
    x"44",
    x"44",
    x"44",
    x"84",
    x"01",
    x"a7",
    x"3e",
    x"ec",
    x"24",
    x"e3",
    x"a4",
    x"81",
    x"10",
    x"23",
    x"0a",
    x"81",
    x"b1",
    x"25",
    x"15",
    x"ec",
    x"a4",
    x"2b",
    x"0d",
    x"20",
    x"04",
    x"ec",
    x"a4",
    x"2a",
    x"07",
    x"43",
    x"53",
    x"c3",
    x"00",
    x"01",
    x"ed",
    x"a4",
    x"ec",
    x"24",
    x"e3",
    x"a4",
    x"ed",
    x"24",
    x"ec",
    x"26",
    x"e3",
    x"22",
    x"81",
    x"07",
    x"23",
    x"0a",
    x"81",
    x"73",
    x"25",
    x"15",
    x"ec",
    x"22",
    x"2b",
    x"0d",
    x"20",
    x"04",
    x"ec",
    x"22",
    x"2a",
    x"07",
    x"43",
    x"53",
    x"c3",
    x"00",
    x"01",
    x"ed",
    x"22",
    x"ec",
    x"26",
    x"e3",
    x"22",
    x"ed",
    x"26",
    x"bd",
    x"d8",
    x"52",
    x"ed",
    x"28",
    x"ce",
    x"3e",
    x"e2",
    x"a6",
    x"3e",
    x"27",
    x"03",
    x"33",
    x"c8",
    x"48",
    x"a6",
    x"26",
    x"84",
    x"03",
    x"c6",
    x"12",
    x"3d",
    x"33",
    x"cb",
    x"ef",
    x"2a",
    x"7e",
    x"d8",
    x"60",
    x"10",
    x"8e",
    x"01",
    x"aa",
    x"9e",
    x"3b",
    x"96",
    x"39",
    x"48",
    x"ae",
    x"86",
    x"30",
    x"02",
    x"39",
    x"bd",
    x"cf",
    x"1d",
    x"8d",
    x"ed",
    x"a6",
    x"84",
    x"27",
    x"f6",
    x"e6",
    x"01",
    x"a1",
    x"24",
    x"10",
    x"26",
    x"00",
    x"b8",
    x"e1",
    x"26",
    x"10",
    x"26",
    x"00",
    x"b2",
    x"ce",
    x"3e",
    x"c0",
    x"a6",
    x"05",
    x"a6",
    x"c6",
    x"94",
    x"52",
    x"27",
    x"dd",
    x"a6",
    x"05",
    x"81",
    x"21",
    x"26",
    x"12",
    x"34",
    x"30",
    x"0c",
    x"3a",
    x"bd",
    x"d1",
    x"4c",
    x"bd",
    x"ce",
    x"cf",
    x"cc",
    x"27",
    x"10",
    x"bd",
    x"db",
    x"0c",
    x"35",
    x"30",
    x"ec",
    x"02",
    x"a7",
    x"24",
    x"e7",
    x"26",
    x"a6",
    x"04",
    x"97",
    x"39",
    x"86",
    x"01",
    x"a7",
    x"3b",
    x"bd",
    x"c5",
    x"25",
    x"bd",
    x"d1",
    x"1a",
    x"7f",
    x"01",
    x"ba",
    x"0f",
    x"32",
    x"7f",
    x"01",
    x"cf",
    x"9e",
    x"3b",
    x"96",
    x"39",
    x"48",
    x"ee",
    x"96",
    x"8e",
    x"1c",
    x"00",
    x"9f",
    x"4e",
    x"17",
    x"00",
    x"f5",
    x"bd",
    x"d2",
    x"4e",
    x"8d",
    x"8c",
    x"10",
    x"8e",
    x"3e",
    x"c0",
    x"a6",
    x"05",
    x"a6",
    x"a6",
    x"94",
    x"52",
    x"27",
    x"02",
    x"8d",
    x"58",
    x"30",
    x"88",
    x"06",
    x"a6",
    x"84",
    x"26",
    x"ef",
    x"8e",
    x"04",
    x"00",
    x"9f",
    x"4e",
    x"17",
    x"00",
    x"e5",
    x"be",
    x"01",
    x"eb",
    x"30",
    x"1c",
    x"de",
    x"53",
    x"bd",
    x"d8",
    x"e2",
    x"96",
    x"39",
    x"27",
    x"17",
    x"8e",
    x"03",
    x"6b",
    x"96",
    x"39",
    x"30",
    x"86",
    x"a6",
    x"84",
    x"94",
    x"52",
    x"26",
    x"0a",
    x"a6",
    x"84",
    x"9a",
    x"52",
    x"a7",
    x"84",
    x"cc",
    x"03",
    x"e8",
    x"8c",
    x"dc",
    x"1b",
    x"bd",
    x"db",
    x"0c",
    x"8e",
    x"04",
    x"55",
    x"ce",
    x"db",
    x"04",
    x"bd",
    x"d8",
    x"e2",
    x"ce",
    x"00",
    x"d0",
    x"86",
    x"24",
    x"d6",
    x"39",
    x"ed",
    x"c4",
    x"bd",
    x"d8",
    x"e2",
    x"7e",
    x"cf",
    x"0f",
    x"30",
    x"88",
    x"06",
    x"7e",
    x"cc",
    x"b6",
    x"39",
    x"34",
    x"50",
    x"ec",
    x"84",
    x"81",
    x"ff",
    x"27",
    x"3e",
    x"c1",
    x"40",
    x"25",
    x"03",
    x"cb",
    x"07",
    x"8c",
    x"c0",
    x"04",
    x"34",
    x"04",
    x"bd",
    x"d8",
    x"56",
    x"1f",
    x"03",
    x"35",
    x"02",
    x"84",
    x"03",
    x"97",
    x"26",
    x"34",
    x"40",
    x"ce",
    x"00",
    x"83",
    x"8e",
    x"df",
    x"0a",
    x"86",
    x"10",
    x"97",
    x"4d",
    x"ec",
    x"81",
    x"ed",
    x"c1",
    x"6f",
    x"c0",
    x"0a",
    x"4d",
    x"26",
    x"f6",
    x"96",
    x"26",
    x"27",
    x"29",
    x"c6",
    x"10",
    x"8d",
    x"0c",
    x"35",
    x"40",
    x"8e",
    x"00",
    x"83",
    x"86",
    x"10",
    x"bd",
    x"d8",
    x"9b",
    x"35",
    x"d0",
    x"8e",
    x"00",
    x"83",
    x"96",
    x"26",
    x"64",
    x"84",
    x"66",
    x"01",
    x"66",
    x"02",
    x"64",
    x"84",
    x"66",
    x"01",
    x"66",
    x"02",
    x"4a",
    x"26",
    x"f1",
    x"30",
    x"03",
    x"5a",
    x"26",
    x"ea",
    x"39",
    x"b6",
    x"ff",
    x"22",
    x"84",
    x"07",
    x"9a",
    x"6a",
    x"b7",
    x"ff",
    x"22",
    x"b7",
    x"ff",
    x"c0",
    x"b7",
    x"ff",
    x"c3",
    x"b7",
    x"ff",
    x"c5",
    x"39",
    x"8e",
    x"ff",
    x"c6",
    x"44",
    x"c6",
    x"07",
    x"44",
    x"25",
    x"03",
    x"a7",
    x"84",
    x"8c",
    x"a7",
    x"01",
    x"30",
    x"02",
    x"5a",
    x"26",
    x"f3",
    x"39",
    x"8e",
    x"1c",
    x"00",
    x"20",
    x"03",
    x"8e",
    x"04",
    x"00",
    x"dc",
    x"1b",
    x"ed",
    x"81",
    x"8c",
    x"34",
    x"00",
    x"26",
    x"f9",
    x"39",
    x"6f",
    x"e2",
    x"8e",
    x"04",
    x"00",
    x"1f",
    x"10",
    x"c5",
    x"1f",
    x"26",
    x"08",
    x"10",
    x"8e",
    x"04",
    x"00",
    x"31",
    x"3f",
    x"26",
    x"fc",
    x"c6",
    x"06",
    x"a6",
    x"89",
    x"18",
    x"00",
    x"a7",
    x"84",
    x"a6",
    x"e4",
    x"26",
    x"05",
    x"86",
    x"55",
    x"a7",
    x"88",
    x"20",
    x"30",
    x"89",
    x"04",
    x"00",
    x"34",
    x"04",
    x"1f",
    x"10",
    x"8a",
    x"02",
    x"b7",
    x"ff",
    x"20",
    x"35",
    x"04",
    x"5a",
    x"26",
    x"df",
    x"30",
    x"89",
    x"e8",
    x"01",
    x"8c",
    x"07",
    x"e0",
    x"25",
    x"04",
    x"86",
    x"ff",
    x"a7",
    x"e4",
    x"8c",
    x"08",
    x"00",
    x"26",
    x"bd",
    x"35",
    x"02",
    x"39",
    x"10",
    x"8e",
    x"01",
    x"aa",
    x"86",
    x"02",
    x"a7",
    x"3b",
    x"86",
    x"10",
    x"a7",
    x"3f",
    x"39",
    x"8e",
    x"ce",
    x"ac",
    x"a6",
    x"80",
    x"2b",
    x"2f",
    x"91",
    x"39",
    x"26",
    x"f8",
    x"10",
    x"8e",
    x"01",
    x"bf",
    x"8e",
    x"01",
    x"ba",
    x"6f",
    x"80",
    x"8c",
    x"01",
    x"cf",
    x"26",
    x"f9",
    x"86",
    x"01",
    x"a7",
    x"3b",
    x"86",
    x"08",
    x"a7",
    x"3f",
    x"cc",
    x"ff",
    x"a8",
    x"ed",
    x"22",
    x"dc",
    x"1b",
    x"ed",
    x"a4",
    x"cc",
    x"74",
    x"65",
    x"a7",
    x"24",
    x"e7",
    x"26",
    x"bd",
    x"d8",
    x"52",
    x"ed",
    x"28",
    x"39",
    x"00",
    x"02",
    x"05",
    x"06",
    x"0a",
    x"0b",
    x"0c",
    x"0d",
    x"0e",
    x"ff",
    x"bd",
    x"ce",
    x"10",
    x"bd",
    x"cd",
    x"e3",
    x"8e",
    x"d2",
    x"5a",
    x"9f",
    x"3b",
    x"0f",
    x"39",
    x"39",
    x"80",
    x"0c",
    x"04",
    x"81",
    x"0a",
    x"89",
    x"0e",
    x"87",
    x"0a",
    x"02",
    x"ff",
    x"c6",
    x"22",
    x"8e",
    x"3e",
    x"c0",
    x"6f",
    x"80",
    x"5a",
    x"26",
    x"fb",
    x"8e",
    x"3e",
    x"c0",
    x"ce",
    x"ce",
    x"ea",
    x"c6",
    x"03",
    x"a6",
    x"c0",
    x"2b",
    x"04",
    x"e7",
    x"86",
    x"20",
    x"f8",
    x"39",
    x"00",
    x"02",
    x"04",
    x"05",
    x"07",
    x"08",
    x"09",
    x"0c",
    x"0d",
    x"0e",
    x"0f",
    x"10",
    x"11",
    x"12",
    x"14",
    x"ff",
    x"10",
    x"8e",
    x"01",
    x"e9",
    x"cc",
    x"02",
    x"14",
    x"bd",
    x"d8",
    x"56",
    x"ed",
    x"22",
    x"86",
    x"07",
    x"a7",
    x"3f",
    x"86",
    x"03",
    x"a7",
    x"3b",
    x"39",
    x"10",
    x"8e",
    x"02",
    x"71",
    x"96",
    x"39",
    x"c6",
    x"19",
    x"3d",
    x"31",
    x"ab",
    x"10",
    x"9f",
    x"3d",
    x"86",
    x"05",
    x"97",
    x"4d",
    x"10",
    x"9e",
    x"3d",
    x"a6",
    x"a4",
    x"94",
    x"52",
    x"27",
    x"12",
    x"bd",
    x"d1",
    x"42",
    x"58",
    x"a6",
    x"21",
    x"3d",
    x"ce",
    x"de",
    x"b3",
    x"33",
    x"cb",
    x"c6",
    x"0a",
    x"d7",
    x"26",
    x"8d",
    x"07",
    x"31",
    x"25",
    x"0a",
    x"4d",
    x"26",
    x"e2",
    x"39",
    x"ec",
    x"c1",
    x"aa",
    x"84",
    x"ea",
    x"01",
    x"ed",
    x"84",
    x"30",
    x"88",
    x"20",
    x"0a",
    x"26",
    x"26",
    x"f1",
    x"39",
    x"10",
    x"8e",
    x"01",
    x"ef",
    x"96",
    x"40",
    x"27",
    x"02",
    x"31",
    x"2d",
    x"03",
    x"40",
    x"a6",
    x"a4",
    x"27",
    x"4a",
    x"2b",
    x"49",
    x"4a",
    x"27",
    x"5c",
    x"ae",
    x"2a",
    x"30",
    x"89",
    x"18",
    x"c0",
    x"a6",
    x"84",
    x"a4",
    x"2c",
    x"bd",
    x"ca",
    x"9b",
    x"26",
    x"4b",
    x"a6",
    x"88",
    x"20",
    x"a4",
    x"2c",
    x"bd",
    x"ca",
    x"9b",
    x"26",
    x"41",
    x"ec",
    x"23",
    x"e3",
    x"21",
    x"ed",
    x"23",
    x"cc",
    x"02",
    x"00",
    x"ed",
    x"21",
    x"a6",
    x"23",
    x"e6",
    x"25",
    x"bd",
    x"d8",
    x"56",
    x"ed",
    x"28",
    x"17",
    x"00",
    x"9d",
    x"ae",
    x"28",
    x"af",
    x"2a",
    x"ee",
    x"26",
    x"c6",
    x"06",
    x"d7",
    x"26",
    x"8d",
    x"9f",
    x"31",
    x"a8",
    x"1a",
    x"10",
    x"8c",
    x"02",
    x"71",
    x"25",
    x"b2",
    x"39",
    x"6a",
    x"a4",
    x"a6",
    x"a4",
    x"84",
    x"02",
    x"27",
    x"05",
    x"cc",
    x"00",
    x"80",
    x"20",
    x"03",
    x"cc",
    x"ff",
    x"80",
    x"ed",
    x"21",
    x"20",
    x"bf",
    x"8d",
    x"71",
    x"c6",
    x"a8",
    x"e7",
    x"a4",
    x"8e",
    x"d0",
    x"5d",
    x"96",
    x"39",
    x"48",
    x"ae",
    x"86",
    x"86",
    x"03",
    x"e6",
    x"80",
    x"bd",
    x"dc",
    x"1f",
    x"3d",
    x"3a",
    x"e6",
    x"84",
    x"bd",
    x"dc",
    x"1f",
    x"86",
    x"08",
    x"3d",
    x"eb",
    x"02",
    x"96",
    x"3a",
    x"81",
    x"03",
    x"25",
    x"02",
    x"c4",
    x"fe",
    x"a6",
    x"01",
    x"a7",
    x"23",
    x"e7",
    x"25",
    x"8b",
    x"06",
    x"cb",
    x"04",
    x"bd",
    x"d8",
    x"56",
    x"1f",
    x"01",
    x"a6",
    x"89",
    x"18",
    x"00",
    x"8e",
    x"d8",
    x"4a",
    x"e6",
    x"25",
    x"c4",
    x"03",
    x"a4",
    x"85",
    x"bd",
    x"c8",
    x"b9",
    x"27",
    x"02",
    x"6a",
    x"25",
    x"a6",
    x"23",
    x"e6",
    x"25",
    x"bd",
    x"d8",
    x"56",
    x"ed",
    x"28",
    x"ed",
    x"2a",
    x"ce",
    x"df",
    x"2a",
    x"a6",
    x"25",
    x"84",
    x"03",
    x"8e",
    x"d0",
    x"31",
    x"e6",
    x"86",
    x"e7",
    x"2c",
    x"c6",
    x"0c",
    x"3d",
    x"33",
    x"cb",
    x"ef",
    x"26",
    x"16",
    x"ff",
    x"7d",
    x"f0",
    x"3c",
    x"0f",
    x"03",
    x"ae",
    x"2a",
    x"ee",
    x"26",
    x"86",
    x"06",
    x"97",
    x"26",
    x"a6",
    x"c0",
    x"43",
    x"a4",
    x"84",
    x"aa",
    x"89",
    x"18",
    x"00",
    x"a7",
    x"84",
    x"e6",
    x"c0",
    x"27",
    x"09",
    x"53",
    x"e4",
    x"01",
    x"ea",
    x"89",
    x"18",
    x"01",
    x"e7",
    x"01",
    x"30",
    x"88",
    x"20",
    x"0a",
    x"26",
    x"26",
    x"e1",
    x"39",
    x"d0",
    x"73",
    x"d0",
    x"89",
    x"d0",
    x"9c",
    x"d0",
    x"ac",
    x"d0",
    x"bf",
    x"d0",
    x"cf",
    x"d0",
    x"df",
    x"d0",
    x"e6",
    x"d0",
    x"fc",
    x"d1",
    x"0c",
    x"d1",
    x"16",
    x"06",
    x"0c",
    x"11",
    x"0f",
    x"09",
    x"3e",
    x"27",
    x"01",
    x"6b",
    x"0f",
    x"05",
    x"6b",
    x"2f",
    x"01",
    x"98",
    x"1f",
    x"01",
    x"98",
    x"3f",
    x"01",
    x"98",
    x"5f",
    x"05",
    x"05",
    x"11",
    x"0f",
    x"04",
    x"11",
    x"4f",
    x"05",
    x"3e",
    x"0f",
    x"01",
    x"3e",
    x"4f",
    x"01",
    x"6b",
    x"67",
    x"02",
    x"98",
    x"47",
    x"04",
    x"0c",
    x"11",
    x"0f",
    x"02",
    x"3e",
    x"0f",
    x"01",
    x"3e",
    x"37",
    x"09",
    x"6b",
    x"27",
    x"04",
    x"98",
    x"0f",
    x"05",
    x"0c",
    x"11",
    x"0f",
    x"03",
    x"3e",
    x"0f",
    x"06",
    x"3e",
    x"3f",
    x"03",
    x"6b",
    x"0f",
    x"00",
    x"98",
    x"0f",
    x"01",
    x"98",
    x"2f",
    x"04",
    x"0c",
    x"11",
    x"0f",
    x"01",
    x"3e",
    x"0f",
    x"08",
    x"4d",
    x"1f",
    x"01",
    x"98",
    x"2f",
    x"01",
    x"98",
    x"57",
    x"04",
    x"0c",
    x"11",
    x"0f",
    x"01",
    x"3e",
    x"67",
    x"0a",
    x"6b",
    x"1f",
    x"01",
    x"98",
    x"0f",
    x"02",
    x"98",
    x"47",
    x"01",
    x"0c",
    x"11",
    x"0f",
    x"09",
    x"5c",
    x"27",
    x"06",
    x"05",
    x"11",
    x"0f",
    x"01",
    x"20",
    x"3f",
    x"04",
    x"11",
    x"4f",
    x"00",
    x"5c",
    x"27",
    x"00",
    x"5c",
    x"57",
    x"00",
    x"6b",
    x"2f",
    x"00",
    x"6b",
    x"4f",
    x"04",
    x"0c",
    x"11",
    x"0f",
    x"08",
    x"3e",
    x"2f",
    x"0a",
    x"5c",
    x"0f",
    x"0a",
    x"7a",
    x"1f",
    x"0a",
    x"98",
    x"0f",
    x"02",
    x"0c",
    x"11",
    x"0f",
    x"03",
    x"3e",
    x"0f",
    x"05",
    x"5c",
    x"37",
    x"00",
    x"0c",
    x"11",
    x"0e",
    x"4f",
    x"c6",
    x"0a",
    x"8d",
    x"18",
    x"96",
    x"3a",
    x"27",
    x"04",
    x"c6",
    x"0a",
    x"20",
    x"09",
    x"d6",
    x"39",
    x"c1",
    x"05",
    x"24",
    x"02",
    x"c6",
    x"05",
    x"5c",
    x"d7",
    x"3f",
    x"86",
    x"01",
    x"8d",
    x"01",
    x"39",
    x"8e",
    x"01",
    x"ef",
    x"a7",
    x"84",
    x"30",
    x"0d",
    x"5a",
    x"26",
    x"f9",
    x"39",
    x"ec",
    x"22",
    x"bd",
    x"d8",
    x"56",
    x"1f",
    x"01",
    x"c6",
    x"0a",
    x"39",
    x"86",
    x"ff",
    x"8e",
    x"02",
    x"71",
    x"c6",
    x"32",
    x"6f",
    x"84",
    x"6f",
    x"01",
    x"a7",
    x"04",
    x"30",
    x"05",
    x"5a",
    x"26",
    x"f5",
    x"8e",
    x"02",
    x"71",
    x"ce",
    x"d1",
    x"c2",
    x"96",
    x"3a",
    x"27",
    x"03",
    x"ce",
    x"d1",
    x"d6",
    x"c6",
    x"0a",
    x"86",
    x"02",
    x"a7",
    x"01",
    x"a7",
    x"06",
    x"a6",
    x"c0",
    x"a7",
    x"04",
    x"a6",
    x"c0",
    x"a7",
    x"09",
    x"30",
    x"88",
    x"19",
    x"5a",
    x"26",
    x"ec",
    x"ce",
    x"d1",
    x"ea",
    x"c6",
    x"0a",
    x"d7",
    x"26",
    x"8e",
    x"02",
    x"71",
    x"c6",
    x"05",
    x"d7",
    x"4d",
    x"34",
    x"10",
    x"d6",
    x"4d",
    x"5a",
    x"86",
    x"05",
    x"3d",
    x"30",
    x"8b",
    x"86",
    x"03",
    x"a7",
    x"84",
    x"d6",
    x"4d",
    x"5a",
    x"1f",
    x"98",
    x"48",
    x"ec",
    x"c6",
    x"ed",
    x"02",
    x"e6",
    x"01",
    x"26",
    x"07",
    x"bd",
    x"dc",
    x"39",
    x"c4",
    x"01",
    x"e7",
    x"01",
    x"35",
    x"10",
    x"0a",
    x"4d",
    x"26",
    x"d7",
    x"30",
    x"88",
    x"19",
    x"33",
    x"4a",
    x"0a",
    x"26",
    x"26",
    x"ca",
    x"39",
    x"01",
    x"03",
    x"1e",
    x"1c",
    x"13",
    x"06",
    x"0b",
    x"0a",
    x"15",
    x"1a",
    x"16",
    x"17",
    x"18",
    x"19",
    x"1b",
    x"21",
    x"1d",
    x"ff",
    x"1f",
    x"20",
    x"01",
    x"03",
    x"1e",
    x"1c",
    x"06",
    x"13",
    x"0a",
    x"0b",
    x"15",
    x"1a",
    x"17",
    x"16",
    x"19",
    x"18",
    x"21",
    x"1b",
    x"1d",
    x"ff",
    x"20",
    x"1f",
    x"3a",
    x"1c",
    x"69",
    x"5c",
    x"65",
    x"20",
    x"91",
    x"30",
    x"91",
    x"50",
    x"23",
    x"34",
    x"23",
    x"48",
    x"38",
    x"64",
    x"97",
    x"3c",
    x"97",
    x"5c",
    x"3a",
    x"60",
    x"44",
    x"1c",
    x"4d",
    x"34",
    x"69",
    x"64",
    x"78",
    x"40",
    x"41",
    x"70",
    x"4b",
    x"24",
    x"6c",
    x"50",
    x"6c",
    x"70",
    x"9d",
    x"0c",
    x"3f",
    x"0c",
    x"6c",
    x"0c",
    x"17",
    x"60",
    x"96",
    x"3c",
    x"96",
    x"64",
    x"14",
    x"6c",
    x"30",
    x"04",
    x"4b",
    x"1c",
    x"5d",
    x"04",
    x"9b",
    x"50",
    x"15",
    x"18",
    x"6a",
    x"6c",
    x"2b",
    x"40",
    x"5f",
    x"18",
    x"93",
    x"34",
    x"30",
    x"0c",
    x"9b",
    x"44",
    x"2c",
    x"3c",
    x"3d",
    x"6c",
    x"9b",
    x"2c",
    x"21",
    x"38",
    x"34",
    x"20",
    x"40",
    x"60",
    x"5d",
    x"1c",
    x"7c",
    x"60",
    x"13",
    x"30",
    x"3d",
    x"38",
    x"44",
    x"18",
    x"96",
    x"38",
    x"96",
    x"60",
    x"86",
    x"01",
    x"97",
    x"20",
    x"cc",
    x"10",
    x"0f",
    x"dd",
    x"21",
    x"7e",
    x"d5",
    x"9e",
    x"d2",
    x"6e",
    x"d2",
    x"7d",
    x"d2",
    x"98",
    x"d2",
    x"bf",
    x"d2",
    x"ec",
    x"d3",
    x"07",
    x"d3",
    x"1c",
    x"d3",
    x"2b",
    x"d3",
    x"3a",
    x"d3",
    x"49",
    x"d3",
    x"5e",
    x"ff",
    x"ff",
    x"a5",
    x"70",
    x"00",
    x"00",
    x"1e",
    x"72",
    x"87",
    x"07",
    x"01",
    x"01",
    x"00",
    x"d3",
    x"a0",
    x"87",
    x"05",
    x"1e",
    x"70",
    x"00",
    x"02",
    x"4b",
    x"72",
    x"a5",
    x"07",
    x"02",
    x"03",
    x"1e",
    x"72",
    x"78",
    x"07",
    x"02",
    x"04",
    x"1e",
    x"05",
    x"78",
    x"70",
    x"06",
    x"1a",
    x"00",
    x"d3",
    x"e4",
    x"a5",
    x"05",
    x"4b",
    x"70",
    x"01",
    x"05",
    x"78",
    x"05",
    x"1e",
    x"70",
    x"01",
    x"06",
    x"78",
    x"72",
    x"78",
    x"07",
    x"03",
    x"07",
    x"4b",
    x"72",
    x"4b",
    x"07",
    x"03",
    x"13",
    x"1e",
    x"72",
    x"1e",
    x"07",
    x"03",
    x"12",
    x"1e",
    x"05",
    x"87",
    x"70",
    x"05",
    x"15",
    x"00",
    x"d4",
    x"26",
    x"78",
    x"05",
    x"78",
    x"70",
    x"02",
    x"08",
    x"a5",
    x"72",
    x"a5",
    x"07",
    x"04",
    x"09",
    x"78",
    x"72",
    x"78",
    x"07",
    x"04",
    x"0a",
    x"4b",
    x"05",
    x"4b",
    x"70",
    x"02",
    x"14",
    x"4b",
    x"72",
    x"4b",
    x"07",
    x"04",
    x"0b",
    x"1e",
    x"05",
    x"1e",
    x"70",
    x"02",
    x"11",
    x"1e",
    x"72",
    x"1e",
    x"07",
    x"04",
    x"10",
    x"00",
    x"d4",
    x"67",
    x"a5",
    x"05",
    x"a5",
    x"70",
    x"03",
    x"0c",
    x"78",
    x"05",
    x"78",
    x"70",
    x"03",
    x"0d",
    x"4b",
    x"05",
    x"4b",
    x"70",
    x"03",
    x"0e",
    x"1e",
    x"05",
    x"1e",
    x"70",
    x"03",
    x"0f",
    x"00",
    x"d4",
    x"a2",
    x"87",
    x"72",
    x"1e",
    x"07",
    x"02",
    x"16",
    x"a5",
    x"05",
    x"3c",
    x"70",
    x"06",
    x"17",
    x"4b",
    x"72",
    x"a5",
    x"07",
    x"07",
    x"1a",
    x"00",
    x"d4",
    x"d9",
    x"78",
    x"72",
    x"1e",
    x"07",
    x"01",
    x"19",
    x"3c",
    x"72",
    x"a5",
    x"07",
    x"05",
    x"18",
    x"00",
    x"d4",
    x"f6",
    x"a5",
    x"05",
    x"4b",
    x"70",
    x"05",
    x"1b",
    x"4b",
    x"72",
    x"a5",
    x"07",
    x"08",
    x"1c",
    x"00",
    x"d5",
    x"2f",
    x"a5",
    x"05",
    x"4b",
    x"70",
    x"07",
    x"1d",
    x"2d",
    x"72",
    x"1e",
    x"07",
    x"09",
    x"1e",
    x"00",
    x"d5",
    x"61",
    x"96",
    x"05",
    x"a5",
    x"70",
    x"08",
    x"20",
    x"1e",
    x"05",
    x"2d",
    x"70",
    x"08",
    x"1f",
    x"a5",
    x"72",
    x"a5",
    x"70",
    x"00",
    x"21",
    x"00",
    x"0f",
    x"80",
    x"06",
    x"0c",
    x"80",
    x"04",
    x"04",
    x"0a",
    x"89",
    x"0b",
    x"03",
    x"80",
    x"08",
    x"0f",
    x"04",
    x"81",
    x"07",
    x"89",
    x"0e",
    x"87",
    x"04",
    x"02",
    x"0f",
    x"19",
    x"19",
    x"17",
    x"01",
    x"0c",
    x"07",
    x"97",
    x"03",
    x"01",
    x"0c",
    x"07",
    x"97",
    x"03",
    x"01",
    x"0c",
    x"07",
    x"09",
    x"98",
    x"03",
    x"09",
    x"98",
    x"03",
    x"09",
    x"18",
    x"1a",
    x"1a",
    x"05",
    x"17",
    x"03",
    x"0d",
    x"80",
    x"03",
    x"0d",
    x"05",
    x"89",
    x"07",
    x"18",
    x"89",
    x"03",
    x"87",
    x"04",
    x"02",
    x"ff",
    x"80",
    x"05",
    x"04",
    x"17",
    x"02",
    x"00",
    x"00",
    x"0d",
    x"00",
    x"04",
    x"0a",
    x"09",
    x"03",
    x"01",
    x"0a",
    x"89",
    x"03",
    x"03",
    x"0f",
    x"04",
    x"81",
    x"04",
    x"89",
    x"0a",
    x"87",
    x"06",
    x"09",
    x"81",
    x"05",
    x"09",
    x"09",
    x"07",
    x"09",
    x"0b",
    x"87",
    x"04",
    x"02",
    x"10",
    x"80",
    x"03",
    x"12",
    x"04",
    x"81",
    x"04",
    x"03",
    x"00",
    x"00",
    x"05",
    x"09",
    x"07",
    x"09",
    x"07",
    x"09",
    x"07",
    x"07",
    x"02",
    x"0d",
    x"07",
    x"09",
    x"09",
    x"07",
    x"18",
    x"01",
    x"89",
    x"07",
    x"0b",
    x"02",
    x"ff",
    x"80",
    x"03",
    x"0c",
    x"80",
    x"04",
    x"0f",
    x"00",
    x"0d",
    x"00",
    x"04",
    x"0a",
    x"09",
    x"03",
    x"01",
    x"0a",
    x"89",
    x"09",
    x"19",
    x"00",
    x"0f",
    x"80",
    x"03",
    x"0c",
    x"00",
    x"00",
    x"04",
    x"0a",
    x"09",
    x"09",
    x"01",
    x"09",
    x"09",
    x"01",
    x"09",
    x"09",
    x"01",
    x"89",
    x"08",
    x"0b",
    x"02",
    x"80",
    x"04",
    x"07",
    x"89",
    x"05",
    x"0b",
    x"87",
    x"03",
    x"02",
    x"0f",
    x"00",
    x"04",
    x"01",
    x"09",
    x"03",
    x"00",
    x"1a",
    x"07",
    x"02",
    x"0c",
    x"05",
    x"89",
    x"08",
    x"0b",
    x"02",
    x"ff",
    x"80",
    x"0c",
    x"04",
    x"0a",
    x"89",
    x"0d",
    x"19",
    x"80",
    x"03",
    x"04",
    x"01",
    x"09",
    x"09",
    x"01",
    x"0f",
    x"04",
    x"01",
    x"01",
    x"00",
    x"87",
    x"05",
    x"02",
    x"12",
    x"00",
    x"0d",
    x"00",
    x"12",
    x"00",
    x"04",
    x"0a",
    x"09",
    x"03",
    x"01",
    x"0a",
    x"09",
    x"03",
    x"01",
    x"0a",
    x"89",
    x"04",
    x"87",
    x"03",
    x"08",
    x"81",
    x"02",
    x"89",
    x"09",
    x"0b",
    x"02",
    x"05",
    x"09",
    x"09",
    x"0b",
    x"02",
    x"00",
    x"07",
    x"09",
    x"09",
    x"0b",
    x"02",
    x"1a",
    x"09",
    x"0b",
    x"02",
    x"ff",
    x"80",
    x"0b",
    x"12",
    x"04",
    x"81",
    x"0a",
    x"89",
    x"0e",
    x"0b",
    x"07",
    x"05",
    x"09",
    x"0b",
    x"07",
    x"05",
    x"09",
    x"0b",
    x"02",
    x"00",
    x"04",
    x"11",
    x"00",
    x"14",
    x"96",
    x"04",
    x"15",
    x"98",
    x"06",
    x"80",
    x"06",
    x"19",
    x"19",
    x"09",
    x"98",
    x"04",
    x"09",
    x"81",
    x"03",
    x"0c",
    x"87",
    x"03",
    x"97",
    x"04",
    x"81",
    x"03",
    x"0c",
    x"87",
    x"03",
    x"1a",
    x"1a",
    x"07",
    x"89",
    x"07",
    x"07",
    x"89",
    x"04",
    x"0b",
    x"02",
    x"ff",
    x"12",
    x"80",
    x"07",
    x"0d",
    x"80",
    x"03",
    x"04",
    x"0a",
    x"89",
    x"03",
    x"03",
    x"00",
    x"04",
    x"0a",
    x"89",
    x"04",
    x"07",
    x"09",
    x"07",
    x"09",
    x"07",
    x"89",
    x"05",
    x"81",
    x"04",
    x"0d",
    x"00",
    x"0f",
    x"80",
    x"07",
    x"04",
    x"01",
    x"0a",
    x"09",
    x"09",
    x"07",
    x"89",
    x"05",
    x"03",
    x"00",
    x"00",
    x"04",
    x"01",
    x"89",
    x"0b",
    x"0b",
    x"02",
    x"00",
    x"07",
    x"09",
    x"09",
    x"87",
    x"07",
    x"02",
    x"ff",
    x"13",
    x"80",
    x"09",
    x"0d",
    x"00",
    x"04",
    x"01",
    x"01",
    x"0a",
    x"89",
    x"0b",
    x"03",
    x"80",
    x"07",
    x"10",
    x"00",
    x"04",
    x"01",
    x"0a",
    x"09",
    x"03",
    x"01",
    x"01",
    x"89",
    x"0e",
    x"87",
    x"0a",
    x"02",
    x"ff",
    x"00",
    x"13",
    x"80",
    x"03",
    x"04",
    x"00",
    x"02",
    x"00",
    x"00",
    x"13",
    x"00",
    x"04",
    x"81",
    x"03",
    x"0a",
    x"09",
    x"03",
    x"81",
    x"05",
    x"89",
    x"07",
    x"07",
    x"07",
    x"05",
    x"07",
    x"02",
    x"02",
    x"07",
    x"07",
    x"09",
    x"01",
    x"09",
    x"01",
    x"09",
    x"09",
    x"07",
    x"09",
    x"07",
    x"09",
    x"01",
    x"01",
    x"84",
    x"03",
    x"08",
    x"01",
    x"01",
    x"89",
    x"06",
    x"87",
    x"06",
    x"05",
    x"09",
    x"0b",
    x"87",
    x"02",
    x"02",
    x"ff",
    x"14",
    x"96",
    x"09",
    x"15",
    x"98",
    x"0b",
    x"0f",
    x"80",
    x"09",
    x"0d",
    x"00",
    x"04",
    x"01",
    x"0a",
    x"89",
    x"09",
    x"86",
    x"07",
    x"0e",
    x"04",
    x"81",
    x"03",
    x"89",
    x"0b",
    x"86",
    x"09",
    x"0e",
    x"04",
    x"81",
    x"03",
    x"89",
    x"0e",
    x"0b",
    x"02",
    x"86",
    x"0a",
    x"89",
    x"0b",
    x"87",
    x"03",
    x"02",
    x"0e",
    x"86",
    x"09",
    x"89",
    x"0b",
    x"87",
    x"04",
    x"02",
    x"ff",
    x"80",
    x"05",
    x"0d",
    x"00",
    x"0d",
    x"00",
    x"0d",
    x"00",
    x"12",
    x"04",
    x"81",
    x"0a",
    x"89",
    x"0a",
    x"9a",
    x"03",
    x"05",
    x"09",
    x"09",
    x"03",
    x"99",
    x"03",
    x"09",
    x"09",
    x"07",
    x"09",
    x"09",
    x"87",
    x"06",
    x"02",
    x"11",
    x"00",
    x"00",
    x"19",
    x"17",
    x"17",
    x"01",
    x"0d",
    x"07",
    x"17",
    x"01",
    x"0d",
    x"07",
    x"17",
    x"01",
    x"0d",
    x"07",
    x"09",
    x"18",
    x"09",
    x"18",
    x"09",
    x"18",
    x"18",
    x"1a",
    x"05",
    x"89",
    x"05",
    x"0b",
    x"02",
    x"ff",
    x"8e",
    x"d5",
    x"bb",
    x"a6",
    x"c0",
    x"2a",
    x"07",
    x"4c",
    x"27",
    x"12",
    x"4a",
    x"e6",
    x"c0",
    x"8c",
    x"c6",
    x"01",
    x"48",
    x"34",
    x"56",
    x"ad",
    x"96",
    x"35",
    x"56",
    x"5a",
    x"26",
    x"f7",
    x"20",
    x"e7",
    x"39",
    x"d5",
    x"f1",
    x"d6",
    x"06",
    x"d6",
    x"20",
    x"d6",
    x"3f",
    x"d6",
    x"4e",
    x"d6",
    x"5e",
    x"d6",
    x"91",
    x"d6",
    x"01",
    x"d6",
    x"2f",
    x"d6",
    x"9b",
    x"d6",
    x"a4",
    x"d6",
    x"ad",
    x"d6",
    x"d4",
    x"d6",
    x"e0",
    x"d6",
    x"ec",
    x"d6",
    x"f8",
    x"d7",
    x"04",
    x"d7",
    x"10",
    x"d7",
    x"1c",
    x"d7",
    x"28",
    x"d6",
    x"6d",
    x"d6",
    x"7f",
    x"d7",
    x"54",
    x"d6",
    x"b6",
    x"d6",
    x"c5",
    x"d6",
    x"ca",
    x"d6",
    x"cf",
    x"ce",
    x"d5",
    x"f7",
    x"7e",
    x"d7",
    x"62",
    x"03",
    x"80",
    x"04",
    x"00",
    x"80",
    x"0a",
    x"03",
    x"80",
    x"07",
    x"00",
    x"ce",
    x"d6",
    x"16",
    x"20",
    x"03",
    x"ce",
    x"d6",
    x"0c",
    x"7e",
    x"d7",
    x"62",
    x"03",
    x"40",
    x"08",
    x"04",
    x"40",
    x"05",
    x"03",
    x"00",
    x"05",
    x"04",
    x"03",
    x"00",
    x"05",
    x"00",
    x"40",
    x"05",
    x"07",
    x"40",
    x"08",
    x"00",
    x"ce",
    x"d6",
    x"25",
    x"20",
    x"0d",
    x"03",
    x"00",
    x"04",
    x"07",
    x"80",
    x"07",
    x"00",
    x"ff",
    x"07",
    x"00",
    x"ce",
    x"d6",
    x"35",
    x"7e",
    x"d7",
    x"62",
    x"03",
    x"ff",
    x"07",
    x"04",
    x"80",
    x"07",
    x"04",
    x"00",
    x"04",
    x"03",
    x"ce",
    x"d6",
    x"44",
    x"20",
    x"0d",
    x"03",
    x"80",
    x"06",
    x"03",
    x"00",
    x"04",
    x"03",
    x"ff",
    x"08",
    x"03",
    x"ce",
    x"d6",
    x"54",
    x"7e",
    x"d7",
    x"62",
    x"03",
    x"80",
    x"06",
    x"03",
    x"ff",
    x"05",
    x"03",
    x"80",
    x"07",
    x"03",
    x"ce",
    x"d6",
    x"63",
    x"20",
    x"ee",
    x"03",
    x"ff",
    x"08",
    x"00",
    x"00",
    x"05",
    x"00",
    x"80",
    x"05",
    x"00",
    x"ce",
    x"d6",
    x"7b",
    x"86",
    x"03",
    x"97",
    x"20",
    x"8d",
    x"1e",
    x"86",
    x"01",
    x"97",
    x"20",
    x"39",
    x"01",
    x"ff",
    x"0a",
    x"03",
    x"ce",
    x"d6",
    x"8d",
    x"86",
    x"03",
    x"97",
    x"20",
    x"8d",
    x"0c",
    x"86",
    x"01",
    x"97",
    x"20",
    x"39",
    x"01",
    x"ff",
    x"0a",
    x"00",
    x"ce",
    x"d6",
    x"97",
    x"7e",
    x"d7",
    x"62",
    x"01",
    x"00",
    x"09",
    x"02",
    x"ce",
    x"d6",
    x"a0",
    x"20",
    x"f4",
    x"01",
    x"00",
    x"09",
    x"06",
    x"ce",
    x"d6",
    x"a9",
    x"20",
    x"eb",
    x"01",
    x"00",
    x"10",
    x"03",
    x"ce",
    x"d6",
    x"b2",
    x"20",
    x"e2",
    x"01",
    x"00",
    x"10",
    x"00",
    x"ce",
    x"d6",
    x"97",
    x"86",
    x"ff",
    x"97",
    x"20",
    x"bd",
    x"d7",
    x"62",
    x"86",
    x"01",
    x"97",
    x"20",
    x"39",
    x"ce",
    x"d6",
    x"a0",
    x"20",
    x"ef",
    x"ce",
    x"d6",
    x"a9",
    x"20",
    x"ea",
    x"ce",
    x"d6",
    x"16",
    x"20",
    x"e5",
    x"8e",
    x"d6",
    x"d9",
    x"20",
    x"5b",
    x"02",
    x"00",
    x"07",
    x"03",
    x"00",
    x"07",
    x"00",
    x"8e",
    x"d6",
    x"e5",
    x"20",
    x"4f",
    x"02",
    x"00",
    x"16",
    x"03",
    x"00",
    x"16",
    x"00",
    x"8e",
    x"d6",
    x"f1",
    x"20",
    x"43",
    x"02",
    x"00",
    x"25",
    x"03",
    x"00",
    x"25",
    x"00",
    x"8e",
    x"d6",
    x"fd",
    x"20",
    x"37",
    x"02",
    x"00",
    x"34",
    x"03",
    x"00",
    x"34",
    x"00",
    x"8e",
    x"d7",
    x"09",
    x"20",
    x"2b",
    x"02",
    x"00",
    x"43",
    x"03",
    x"00",
    x"43",
    x"00",
    x"8e",
    x"d7",
    x"15",
    x"20",
    x"1f",
    x"02",
    x"00",
    x"52",
    x"03",
    x"00",
    x"52",
    x"00",
    x"8e",
    x"d7",
    x"21",
    x"20",
    x"13",
    x"02",
    x"00",
    x"61",
    x"03",
    x"00",
    x"61",
    x"00",
    x"8e",
    x"d7",
    x"2d",
    x"20",
    x"07",
    x"02",
    x"00",
    x"8e",
    x"03",
    x"00",
    x"8e",
    x"00",
    x"34",
    x"10",
    x"ce",
    x"d7",
    x"4c",
    x"8d",
    x"27",
    x"86",
    x"03",
    x"97",
    x"20",
    x"35",
    x"40",
    x"8d",
    x"1f",
    x"ce",
    x"d7",
    x"50",
    x"86",
    x"01",
    x"97",
    x"20",
    x"20",
    x"16",
    x"01",
    x"ff",
    x"06",
    x"03",
    x"01",
    x"ff",
    x"06",
    x"00",
    x"ce",
    x"d6",
    x"97",
    x"86",
    x"03",
    x"97",
    x"20",
    x"8d",
    x"05",
    x"86",
    x"01",
    x"97",
    x"20",
    x"39",
    x"a6",
    x"c0",
    x"97",
    x"24",
    x"0f",
    x"1e",
    x"a6",
    x"c0",
    x"97",
    x"1f",
    x"a6",
    x"c0",
    x"97",
    x"1d",
    x"a6",
    x"c0",
    x"48",
    x"8e",
    x"d7",
    x"7d",
    x"ad",
    x"96",
    x"0a",
    x"24",
    x"26",
    x"ec",
    x"39",
    x"d7",
    x"8d",
    x"d7",
    x"94",
    x"d7",
    x"9d",
    x"d7",
    x"a4",
    x"d7",
    x"ab",
    x"d7",
    x"b4",
    x"d7",
    x"bb",
    x"d7",
    x"c4",
    x"8e",
    x"d7",
    x"ff",
    x"0f",
    x"25",
    x"20",
    x"52",
    x"8e",
    x"d8",
    x"04",
    x"86",
    x"ff",
    x"97",
    x"25",
    x"20",
    x"30",
    x"8e",
    x"d8",
    x"09",
    x"0f",
    x"25",
    x"20",
    x"29",
    x"8e",
    x"d8",
    x"0e",
    x"0f",
    x"25",
    x"20",
    x"3b",
    x"8e",
    x"d8",
    x"13",
    x"86",
    x"ff",
    x"97",
    x"25",
    x"20",
    x"32",
    x"8e",
    x"d8",
    x"18",
    x"0f",
    x"25",
    x"20",
    x"12",
    x"8e",
    x"d8",
    x"1d",
    x"86",
    x"ff",
    x"97",
    x"25",
    x"20",
    x"09",
    x"8e",
    x"d8",
    x"22",
    x"86",
    x"ff",
    x"97",
    x"25",
    x"20",
    x"19",
    x"96",
    x"21",
    x"d6",
    x"1d",
    x"27",
    x"12",
    x"d6",
    x"25",
    x"34",
    x"56",
    x"8d",
    x"4e",
    x"35",
    x"56",
    x"0a",
    x"1d",
    x"27",
    x"06",
    x"ad",
    x"84",
    x"97",
    x"21",
    x"20",
    x"f0",
    x"39",
    x"96",
    x"22",
    x"d6",
    x"1d",
    x"27",
    x"12",
    x"d6",
    x"25",
    x"34",
    x"56",
    x"8d",
    x"35",
    x"35",
    x"56",
    x"0a",
    x"1d",
    x"27",
    x"06",
    x"ad",
    x"84",
    x"97",
    x"22",
    x"20",
    x"f0",
    x"39",
    x"0a",
    x"21",
    x"d3",
    x"1e",
    x"39",
    x"0c",
    x"22",
    x"93",
    x"1e",
    x"39",
    x"0c",
    x"22",
    x"d3",
    x"1e",
    x"39",
    x"0c",
    x"21",
    x"d3",
    x"1e",
    x"39",
    x"0c",
    x"21",
    x"93",
    x"1e",
    x"39",
    x"0a",
    x"22",
    x"d3",
    x"1e",
    x"39",
    x"0a",
    x"22",
    x"93",
    x"1e",
    x"39",
    x"0a",
    x"21",
    x"93",
    x"1e",
    x"39",
    x"dc",
    x"21",
    x"8d",
    x"2b",
    x"1f",
    x"02",
    x"d6",
    x"22",
    x"c4",
    x"03",
    x"ce",
    x"d8",
    x"4a",
    x"30",
    x"44",
    x"96",
    x"20",
    x"2b",
    x"0f",
    x"a6",
    x"86",
    x"a4",
    x"c5",
    x"a7",
    x"e2",
    x"a6",
    x"c5",
    x"43",
    x"a4",
    x"a4",
    x"aa",
    x"e0",
    x"a7",
    x"a4",
    x"39",
    x"c0",
    x"30",
    x"0c",
    x"03",
    x"00",
    x"55",
    x"aa",
    x"ff",
    x"a6",
    x"24",
    x"e6",
    x"26",
    x"58",
    x"44",
    x"56",
    x"44",
    x"56",
    x"44",
    x"56",
    x"d3",
    x"4e",
    x"39",
    x"a6",
    x"3b",
    x"27",
    x"4e",
    x"2b",
    x"4d",
    x"4a",
    x"27",
    x"03",
    x"8d",
    x"4a",
    x"8c",
    x"6c",
    x"3b",
    x"10",
    x"8c",
    x"01",
    x"aa",
    x"26",
    x"1d",
    x"a6",
    x"35",
    x"27",
    x"19",
    x"e6",
    x"26",
    x"cb",
    x"03",
    x"a6",
    x"24",
    x"dd",
    x"21",
    x"0f",
    x"20",
    x"dc",
    x"1b",
    x"dd",
    x"1e",
    x"86",
    x"0c",
    x"97",
    x"1d",
    x"bd",
    x"d7",
    x"a4",
    x"10",
    x"8e",
    x"01",
    x"aa",
    x"ee",
    x"28",
    x"ef",
    x"2c",
    x"ae",
    x"2a",
    x"af",
    x"2e",
    x"a6",
    x"3f",
    x"97",
    x"26",
    x"ec",
    x"c4",
    x"aa",
    x"80",
    x"ea",
    x"80",
    x"ed",
    x"c4",
    x"a6",
    x"42",
    x"aa",
    x"80",
    x"a7",
    x"42",
    x"33",
    x"c8",
    x"20",
    x"0a",
    x"26",
    x"26",
    x"eb",
    x"39",
    x"6f",
    x"3b",
    x"ee",
    x"2c",
    x"ae",
    x"2e",
    x"a6",
    x"3f",
    x"97",
    x"26",
    x"ec",
    x"81",
    x"43",
    x"a4",
    x"c4",
    x"aa",
    x"c9",
    x"18",
    x"00",
    x"53",
    x"e4",
    x"41",
    x"ea",
    x"c9",
    x"18",
    x"01",
    x"ed",
    x"c4",
    x"a6",
    x"80",
    x"43",
    x"a4",
    x"42",
    x"aa",
    x"c9",
    x"18",
    x"02",
    x"a7",
    x"42",
    x"33",
    x"c8",
    x"20",
    x"0a",
    x"26",
    x"26",
    x"dc",
    x"39",
    x"10",
    x"8e",
    x"d9",
    x"08",
    x"c6",
    x"07",
    x"a6",
    x"c0",
    x"2b",
    x"1b",
    x"3d",
    x"31",
    x"ab",
    x"c6",
    x"07",
    x"a6",
    x"a0",
    x"94",
    x"69",
    x"aa",
    x"89",
    x"18",
    x"00",
    x"a7",
    x"84",
    x"30",
    x"88",
    x"20",
    x"5a",
    x"26",
    x"f0",
    x"30",
    x"89",
    x"ff",
    x"21",
    x"20",
    x"db",
    x"39",
    x"30",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"30",
    x"30",
    x"f0",
    x"30",
    x"30",
    x"30",
    x"30",
    x"fc",
    x"30",
    x"cc",
    x"0c",
    x"30",
    x"30",
    x"c0",
    x"fc",
    x"30",
    x"cc",
    x"0c",
    x"3c",
    x"0c",
    x"cc",
    x"30",
    x"0c",
    x"3c",
    x"cc",
    x"fc",
    x"0c",
    x"0c",
    x"0c",
    x"fc",
    x"c0",
    x"c0",
    x"fc",
    x"0c",
    x"cc",
    x"30",
    x"30",
    x"cc",
    x"c0",
    x"f0",
    x"cc",
    x"cc",
    x"30",
    x"fc",
    x"0c",
    x"30",
    x"30",
    x"30",
    x"c0",
    x"c0",
    x"30",
    x"cc",
    x"cc",
    x"30",
    x"cc",
    x"cc",
    x"30",
    x"30",
    x"cc",
    x"cc",
    x"3c",
    x"0c",
    x"cc",
    x"30",
    x"30",
    x"cc",
    x"cc",
    x"fc",
    x"cc",
    x"cc",
    x"cc",
    x"f0",
    x"cc",
    x"cc",
    x"f0",
    x"cc",
    x"cc",
    x"f0",
    x"30",
    x"cc",
    x"c0",
    x"c0",
    x"c0",
    x"cc",
    x"30",
    x"f0",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"f0",
    x"fc",
    x"c0",
    x"c0",
    x"f0",
    x"c0",
    x"c0",
    x"fc",
    x"fc",
    x"c0",
    x"c0",
    x"f0",
    x"c0",
    x"c0",
    x"c0",
    x"30",
    x"cc",
    x"c0",
    x"3c",
    x"cc",
    x"cc",
    x"30",
    x"cc",
    x"cc",
    x"cc",
    x"fc",
    x"cc",
    x"cc",
    x"cc",
    x"fc",
    x"30",
    x"30",
    x"30",
    x"30",
    x"30",
    x"fc",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"0c",
    x"cc",
    x"30",
    x"cc",
    x"cc",
    x"f0",
    x"c0",
    x"f0",
    x"cc",
    x"cc",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"c0",
    x"fc",
    x"cc",
    x"fc",
    x"fc",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"f0",
    x"fc",
    x"fc",
    x"cc",
    x"cc",
    x"30",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"30",
    x"f0",
    x"cc",
    x"cc",
    x"f0",
    x"c0",
    x"c0",
    x"c0",
    x"30",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"fc",
    x"3c",
    x"f0",
    x"cc",
    x"cc",
    x"f0",
    x"f0",
    x"cc",
    x"cc",
    x"30",
    x"cc",
    x"c0",
    x"30",
    x"0c",
    x"cc",
    x"30",
    x"fc",
    x"30",
    x"30",
    x"30",
    x"30",
    x"30",
    x"30",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"30",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"30",
    x"30",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"fc",
    x"fc",
    x"cc",
    x"cc",
    x"cc",
    x"30",
    x"30",
    x"30",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"cc",
    x"30",
    x"30",
    x"30",
    x"30",
    x"fc",
    x"0c",
    x"30",
    x"30",
    x"30",
    x"c0",
    x"fc",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"c0",
    x"c0",
    x"00",
    x"c0",
    x"c0",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"30",
    x"30",
    x"0d",
    x"18",
    x"20",
    x"17",
    x"15",
    x"0a",
    x"17",
    x"0d",
    x"24",
    x"1f",
    x"01",
    x"26",
    x"01",
    x"ff",
    x"20",
    x"1b",
    x"12",
    x"1d",
    x"1d",
    x"0e",
    x"17",
    x"24",
    x"0b",
    x"22",
    x"25",
    x"ff",
    x"16",
    x"12",
    x"0c",
    x"11",
    x"0a",
    x"0e",
    x"15",
    x"24",
    x"0a",
    x"12",
    x"0c",
    x"11",
    x"15",
    x"16",
    x"0a",
    x"22",
    x"1b",
    x"ff",
    x"0c",
    x"18",
    x"19",
    x"22",
    x"1b",
    x"12",
    x"10",
    x"11",
    x"1d",
    x"24",
    x"01",
    x"09",
    x"08",
    x"03",
    x"ff",
    x"1c",
    x"19",
    x"0e",
    x"0c",
    x"1d",
    x"1b",
    x"0a",
    x"15",
    x"24",
    x"0a",
    x"1c",
    x"1c",
    x"18",
    x"0c",
    x"12",
    x"0a",
    x"1d",
    x"0e",
    x"1c",
    x"ff",
    x"15",
    x"12",
    x"0c",
    x"0e",
    x"17",
    x"1c",
    x"0e",
    x"0d",
    x"24",
    x"1d",
    x"18",
    x"24",
    x"ff",
    x"1d",
    x"0a",
    x"17",
    x"0d",
    x"22",
    x"24",
    x"0c",
    x"18",
    x"1b",
    x"19",
    x"18",
    x"1b",
    x"0a",
    x"1d",
    x"12",
    x"18",
    x"17",
    x"ff",
    x"0a",
    x"15",
    x"15",
    x"24",
    x"1b",
    x"12",
    x"10",
    x"11",
    x"1d",
    x"1c",
    x"24",
    x"1b",
    x"0e",
    x"1c",
    x"0e",
    x"1b",
    x"1f",
    x"0e",
    x"0d",
    x"ff",
    x"18",
    x"17",
    x"0e",
    x"24",
    x"19",
    x"15",
    x"0a",
    x"22",
    x"0e",
    x"1b",
    x"ff",
    x"1d",
    x"20",
    x"18",
    x"24",
    x"19",
    x"15",
    x"0a",
    x"22",
    x"0e",
    x"1b",
    x"ff",
    x"11",
    x"12",
    x"10",
    x"11",
    x"24",
    x"1c",
    x"0c",
    x"18",
    x"1b",
    x"0e",
    x"ff",
    x"19",
    x"15",
    x"0a",
    x"22",
    x"0e",
    x"1b",
    x"24",
    x"18",
    x"17",
    x"0e",
    x"ff",
    x"19",
    x"15",
    x"0a",
    x"22",
    x"0e",
    x"1b",
    x"24",
    x"1d",
    x"20",
    x"18",
    x"ff",
    x"19",
    x"15",
    x"01",
    x"ff",
    x"19",
    x"15",
    x"02",
    x"ff",
    x"10",
    x"0e",
    x"1d",
    x"24",
    x"1b",
    x"0e",
    x"0a",
    x"0d",
    x"22",
    x"24",
    x"19",
    x"15",
    x"0a",
    x"22",
    x"0e",
    x"1b",
    x"24",
    x"18",
    x"17",
    x"0e",
    x"ff",
    x"10",
    x"0e",
    x"1d",
    x"24",
    x"1b",
    x"0e",
    x"0a",
    x"0d",
    x"22",
    x"24",
    x"19",
    x"15",
    x"0a",
    x"22",
    x"0e",
    x"1b",
    x"24",
    x"1d",
    x"20",
    x"18",
    x"ff",
    x"0c",
    x"11",
    x"0a",
    x"16",
    x"0b",
    x"0e",
    x"1b",
    x"ff",
    x"8d",
    x"47",
    x"ce",
    x"db",
    x"32",
    x"96",
    x"52",
    x"84",
    x"02",
    x"ee",
    x"c6",
    x"8d",
    x"79",
    x"8e",
    x"1b",
    x"03",
    x"8d",
    x"03",
    x"7e",
    x"d8",
    x"e2",
    x"a6",
    x"c4",
    x"2b",
    x"08",
    x"26",
    x"0a",
    x"33",
    x"41",
    x"30",
    x"01",
    x"20",
    x"f4",
    x"33",
    x"5f",
    x"30",
    x"1f",
    x"39",
    x"00",
    x"bb",
    x"00",
    x"c3",
    x"34",
    x"10",
    x"8d",
    x"1b",
    x"35",
    x"10",
    x"ce",
    x"00",
    x"cb",
    x"8d",
    x"03",
    x"7e",
    x"d8",
    x"e2",
    x"1f",
    x"32",
    x"a6",
    x"a0",
    x"2b",
    x"08",
    x"26",
    x"08",
    x"86",
    x"24",
    x"a7",
    x"3f",
    x"20",
    x"f4",
    x"6f",
    x"3e",
    x"39",
    x"dd",
    x"6e",
    x"c6",
    x"07",
    x"8e",
    x"00",
    x"cb",
    x"6f",
    x"80",
    x"5a",
    x"26",
    x"fb",
    x"8e",
    x"00",
    x"cd",
    x"cc",
    x"27",
    x"10",
    x"8d",
    x"14",
    x"cc",
    x"03",
    x"e8",
    x"8d",
    x"0f",
    x"cc",
    x"00",
    x"64",
    x"8d",
    x"0a",
    x"cc",
    x"00",
    x"0a",
    x"8d",
    x"05",
    x"d6",
    x"6f",
    x"e7",
    x"84",
    x"39",
    x"0f",
    x"6b",
    x"dd",
    x"6c",
    x"dc",
    x"6e",
    x"dd",
    x"6e",
    x"93",
    x"6c",
    x"25",
    x"04",
    x"0c",
    x"6b",
    x"20",
    x"f6",
    x"96",
    x"6b",
    x"a7",
    x"80",
    x"39",
    x"5f",
    x"8e",
    x"00",
    x"d2",
    x"33",
    x"47",
    x"a6",
    x"c2",
    x"cb",
    x"f0",
    x"a9",
    x"82",
    x"19",
    x"1f",
    x"89",
    x"84",
    x"0f",
    x"a7",
    x"c4",
    x"8c",
    x"00",
    x"cb",
    x"26",
    x"ee",
    x"cb",
    x"f0",
    x"39",
    x"ce",
    x"db",
    x"c1",
    x"ec",
    x"c1",
    x"2b",
    x"0c",
    x"ae",
    x"c1",
    x"10",
    x"ae",
    x"c1",
    x"8d",
    x"1f",
    x"4a",
    x"26",
    x"fb",
    x"20",
    x"f0",
    x"39",
    x"0a",
    x"10",
    x"dc",
    x"d7",
    x"34",
    x"00",
    x"0a",
    x"05",
    x"de",
    x"17",
    x"3b",
    x"80",
    x"02",
    x"08",
    x"de",
    x"7b",
    x"3d",
    x"d8",
    x"02",
    x"06",
    x"de",
    x"9b",
    x"3e",
    x"e2",
    x"ff",
    x"34",
    x"46",
    x"4f",
    x"ed",
    x"e3",
    x"34",
    x"16",
    x"6f",
    x"22",
    x"ec",
    x"81",
    x"6d",
    x"64",
    x"27",
    x"0c",
    x"44",
    x"56",
    x"66",
    x"22",
    x"44",
    x"56",
    x"66",
    x"22",
    x"6a",
    x"64",
    x"20",
    x"f0",
    x"ed",
    x"a4",
    x"31",
    x"23",
    x"a6",
    x"e4",
    x"a7",
    x"64",
    x"6a",
    x"65",
    x"26",
    x"e0",
    x"35",
    x"56",
    x"4c",
    x"81",
    x"04",
    x"26",
    x"d5",
    x"58",
    x"3a",
    x"35",
    x"c6",
    x"35",
    x"10",
    x"96",
    x"50",
    x"84",
    x"02",
    x"10",
    x"27",
    x"e4",
    x"55",
    x"0a",
    x"50",
    x"1f",
    x"20",
    x"34",
    x"16",
    x"7e",
    x"c6",
    x"10",
    x"34",
    x"12",
    x"4f",
    x"dd",
    x"64",
    x"43",
    x"59",
    x"25",
    x"05",
    x"43",
    x"06",
    x"64",
    x"20",
    x"f8",
    x"03",
    x"64",
    x"8d",
    x"08",
    x"d4",
    x"64",
    x"d1",
    x"65",
    x"22",
    x"f8",
    x"35",
    x"92",
    x"34",
    x"10",
    x"9e",
    x"61",
    x"30",
    x"01",
    x"8c",
    x"df",
    x"5a",
    x"25",
    x"03",
    x"8e",
    x"c0",
    x"00",
    x"9f",
    x"61",
    x"e6",
    x"84",
    x"35",
    x"90",
    x"b6",
    x"ff",
    x"02",
    x"0c",
    x"14",
    x"0c",
    x"63",
    x"3b",
    x"ce",
    x"ff",
    x"01",
    x"8d",
    x"00",
    x"a6",
    x"c4",
    x"84",
    x"f7",
    x"54",
    x"24",
    x"02",
    x"8a",
    x"08",
    x"a7",
    x"c1",
    x"39",
    x"8d",
    x"66",
    x"8e",
    x"00",
    x"14",
    x"c6",
    x"01",
    x"d7",
    x"10",
    x"96",
    x"52",
    x"84",
    x"02",
    x"34",
    x"02",
    x"eb",
    x"e0",
    x"8d",
    x"dc",
    x"cc",
    x"40",
    x"80",
    x"97",
    x"11",
    x"ca",
    x"02",
    x"f7",
    x"ff",
    x"20",
    x"c8",
    x"02",
    x"b6",
    x"ff",
    x"00",
    x"2b",
    x"03",
    x"d0",
    x"11",
    x"8c",
    x"db",
    x"11",
    x"96",
    x"11",
    x"44",
    x"81",
    x"01",
    x"26",
    x"e6",
    x"e7",
    x"82",
    x"d6",
    x"10",
    x"5a",
    x"2a",
    x"d0",
    x"ec",
    x"84",
    x"0f",
    x"15",
    x"54",
    x"54",
    x"27",
    x"07",
    x"c1",
    x"3f",
    x"26",
    x"07",
    x"c6",
    x"03",
    x"8c",
    x"c6",
    x"01",
    x"d7",
    x"15",
    x"44",
    x"44",
    x"27",
    x"07",
    x"81",
    x"3f",
    x"26",
    x"07",
    x"86",
    x"02",
    x"8c",
    x"86",
    x"04",
    x"97",
    x"15",
    x"86",
    x"02",
    x"b7",
    x"ff",
    x"20",
    x"5f",
    x"8d",
    x"8e",
    x"b6",
    x"ff",
    x"23",
    x"8a",
    x"08",
    x"20",
    x"05",
    x"b6",
    x"ff",
    x"23",
    x"84",
    x"f7",
    x"b7",
    x"ff",
    x"23",
    x"39",
    x"0a",
    x"80",
    x"2a",
    x"a0",
    x"15",
    x"c0",
    x"2d",
    x"a0",
    x"2d",
    x"d0",
    x"17",
    x"a0",
    x"0f",
    x"e0",
    x"1a",
    x"80",
    x"1a",
    x"c0",
    x"1a",
    x"80",
    x"1f",
    x"80",
    x"0f",
    x"80",
    x"0a",
    x"c0",
    x"0a",
    x"80",
    x"0f",
    x"c0",
    x"0f",
    x"e0",
    x"0a",
    x"80",
    x"2a",
    x"a0",
    x"15",
    x"c0",
    x"2d",
    x"a0",
    x"2d",
    x"d0",
    x"17",
    x"a0",
    x"0f",
    x"e0",
    x"0a",
    x"80",
    x"3a",
    x"d8",
    x"7a",
    x"f8",
    x"6a",
    x"f8",
    x"0a",
    x"a8",
    x"0a",
    x"a8",
    x"2a",
    x"38",
    x"6a",
    x"38",
    x"60",
    x"00",
    x"00",
    x"00",
    x"0a",
    x"80",
    x"2a",
    x"a0",
    x"15",
    x"c0",
    x"2d",
    x"a0",
    x"2d",
    x"d0",
    x"17",
    x"a0",
    x"0f",
    x"e6",
    x"fa",
    x"fe",
    x"fa",
    x"fe",
    x"0a",
    x"a0",
    x"0a",
    x"aa",
    x"3a",
    x"ae",
    x"6a",
    x"0e",
    x"60",
    x"00",
    x"00",
    x"00",
    x"0a",
    x"80",
    x"2a",
    x"a0",
    x"15",
    x"c0",
    x"2d",
    x"a0",
    x"2d",
    x"d0",
    x"17",
    x"a0",
    x"0f",
    x"e0",
    x"0a",
    x"80",
    x"7a",
    x"d8",
    x"7a",
    x"f8",
    x"6a",
    x"f0",
    x"0a",
    x"a0",
    x"6a",
    x"a0",
    x"68",
    x"50",
    x"60",
    x"70",
    x"00",
    x"38",
    x"0a",
    x"c0",
    x"1a",
    x"b0",
    x"15",
    x"58",
    x"35",
    x"58",
    x"35",
    x"58",
    x"15",
    x"58",
    x"35",
    x"b8",
    x"6a",
    x"b0",
    x"ea",
    x"a0",
    x"6a",
    x"a0",
    x"2a",
    x"a0",
    x"2a",
    x"a0",
    x"28",
    x"a0",
    x"1c",
    x"a0",
    x"00",
    x"a0",
    x"01",
    x"c0",
    x"1a",
    x"80",
    x"6a",
    x"c0",
    x"d5",
    x"40",
    x"d5",
    x"60",
    x"d5",
    x"60",
    x"d5",
    x"40",
    x"ea",
    x"e0",
    x"6a",
    x"b0",
    x"2a",
    x"b8",
    x"2a",
    x"b0",
    x"2a",
    x"a0",
    x"2a",
    x"a0",
    x"28",
    x"a0",
    x"29",
    x"c0",
    x"28",
    x"00",
    x"1c",
    x"00",
    x"02",
    x"a0",
    x"0a",
    x"a8",
    x"07",
    x"50",
    x"0b",
    x"68",
    x"17",
    x"68",
    x"0b",
    x"d0",
    x"0f",
    x"e0",
    x"02",
    x"b0",
    x"06",
    x"b0",
    x"02",
    x"b0",
    x"03",
    x"f0",
    x"03",
    x"e0",
    x"06",
    x"a0",
    x"02",
    x"a0",
    x"07",
    x"e0",
    x"0f",
    x"e0",
    x"02",
    x"a0",
    x"0a",
    x"a8",
    x"07",
    x"50",
    x"0b",
    x"68",
    x"17",
    x"68",
    x"0b",
    x"d0",
    x"0f",
    x"f0",
    x"02",
    x"a0",
    x"1a",
    x"bc",
    x"1e",
    x"b7",
    x"1e",
    x"a6",
    x"0a",
    x"a0",
    x"0a",
    x"a0",
    x"1c",
    x"ae",
    x"1c",
    x"ae",
    x"00",
    x"06",
    x"00",
    x"00",
    x"02",
    x"a0",
    x"0a",
    x"a8",
    x"07",
    x"50",
    x"0b",
    x"68",
    x"17",
    x"68",
    x"0b",
    x"d0",
    x"6f",
    x"e0",
    x"7e",
    x"bf",
    x"7e",
    x"bf",
    x"0a",
    x"a0",
    x"6a",
    x"a0",
    x"7a",
    x"ae",
    x"78",
    x"ae",
    x"00",
    x"06",
    x"00",
    x"00",
    x"02",
    x"a0",
    x"0a",
    x"a8",
    x"07",
    x"50",
    x"0b",
    x"68",
    x"17",
    x"68",
    x"0b",
    x"d0",
    x"0f",
    x"e0",
    x"02",
    x"a0",
    x"1a",
    x"be",
    x"1e",
    x"be",
    x"1e",
    x"a6",
    x"0a",
    x"a0",
    x"0a",
    x"ae",
    x"08",
    x"ae",
    x"1c",
    x"06",
    x"1c",
    x"00",
    x"3f",
    x"f0",
    x"3f",
    x"f0",
    x"3f",
    x"c0",
    x"3f",
    x"c0",
    x"0f",
    x"c0",
    x"3f",
    x"f0",
    x"3f",
    x"f0",
    x"0f",
    x"c0",
    x"6f",
    x"f8",
    x"3f",
    x"38",
    x"0f",
    x"c0",
    x"3f",
    x"f0",
    x"0f",
    x"f6",
    x"0f",
    x"f0",
    x"7f",
    x"0e",
    x"3f",
    x"f0",
    x"3f",
    x"f0",
    x"0f",
    x"c0",
    x"6f",
    x"f0",
    x"6c",
    x"70",
    x"3f",
    x"f0",
    x"3f",
    x"fc",
    x"ff",
    x"f0",
    x"3f",
    x"f0",
    x"3c",
    x"f0",
    x"ff",
    x"c0",
    x"ff",
    x"f0",
    x"ff",
    x"f0",
    x"3f",
    x"f0",
    x"3f",
    x"c0",
    x"0f",
    x"fc",
    x"1f",
    x"f8",
    x"03",
    x"f0",
    x"03",
    x"f0",
    x"03",
    x"f0",
    x"0f",
    x"f8",
    x"1f",
    x"f8",
    x"03",
    x"f0",
    x"1f",
    x"f6",
    x"1c",
    x"fe",
    x"03",
    x"f0",
    x"0f",
    x"f8",
    x"6f",
    x"f0",
    x"0f",
    x"f0",
    x"7c",
    x"fe",
    x"0f",
    x"f8",
    x"1f",
    x"f8",
    x"03",
    x"f0",
    x"1f",
    x"f6",
    x"0c",
    x"fe",
    x"01",
    x"00",
    x"05",
    x"40",
    x"0d",
    x"60",
    x"15",
    x"50",
    x"15",
    x"50",
    x"0d",
    x"60",
    x"05",
    x"40",
    x"01",
    x"00",
    x"00",
    x"00",
    x"00",
    x"00",
    x"05",
    x"40",
    x"35",
    x"58",
    x"55",
    x"54",
    x"55",
    x"54",
    x"35",
    x"58",
    x"05",
    x"40",
    x"c1",
    x"83",
    x"f3",
    x"cf",
    x"3f",
    x"fc",
    x"0f",
    x"f0",
    x"03",
    x"c0",
    x"01",
    x"80",
    x"01",
    x"80",
    x"03",
    x"c0",
    x"0f",
    x"f0",
    x"3f",
    x"fc",
    x"f3",
    x"cf",
    x"c1",
    x"83",
    x"11",
    x"10",
    x"1e",
    x"e4",
    x"0a",
    x"d8",
    x"07",
    x"f0",
    x"0d",
    x"6c",
    x"1a",
    x"b2",
    x"3a",
    x"b8",
    x"3a",
    x"b8",
    x"3a",
    x"b8",
    x"1f",
    x"f0",
    x"02",
    x"80",
    x"2a",
    x"a8",
    x"aa",
    x"aa",
    x"aa",
    x"aa",
    x"2a",
    x"a8",
    x"2a",
    x"a8",
    x"0a",
    x"a0",
    x"0a",
    x"a0",
    x"02",
    x"80",
    x"02",
    x"80",
    x"00",
    x"00",
    x"20",
    x"00",
    x"28",
    x"00",
    x"88",
    x"00",
    x"8b",
    x"55",
    x"8a",
    x"aa",
    x"8b",
    x"55",
    x"88",
    x"33",
    x"28",
    x"33",
    x"20",
    x"00",
    x"04",
    x"00",
    x"00",
    x"03",
    x"07",
    x"00",
    x"31",
    x"06",
    x"00",
    x"18",
    x"04",
    x"c0",
    x"09",
    x"50",
    x"80",
    x"05",
    x"54",
    x"00",
    x"16",
    x"5c",
    x"00",
    x"39",
    x"55",
    x"00",
    x"da",
    x"ab",
    x"c0",
    x"2a",
    x"80",
    x"aa",
    x"a0",
    x"af",
    x"a0",
    x"b5",
    x"e0",
    x"af",
    x"a0",
    x"aa",
    x"a0",
    x"a5",
    x"a0",
    x"9a",
    x"60",
    x"9a",
    x"60",
    x"a5",
    x"a0",
    x"aa",
    x"a0",
    x"aa",
    x"a0",
    x"aa",
    x"a0",
    x"aa",
    x"a0",
    x"aa",
    x"a0",
    x"aa",
    x"a0",
    x"00",
    x"00",
    x"40",
    x"00",
    x"60",
    x"00",
    x"f0",
    x"00",
    x"f0",
    x"00",
    x"60",
    x"00",
    x"00",
    x"00",
    x"10",
    x"00",
    x"18",
    x"00",
    x"3c",
    x"00",
    x"3c",
    x"00",
    x"18",
    x"00",
    x"00",
    x"00",
    x"04",
    x"00",
    x"06",
    x"00",
    x"0f",
    x"00",
    x"0f",
    x"00",
    x"06",
    x"00",
    x"00",
    x"00",
    x"01",
    x"00",
    x"01",
    x"80",
    x"03",
    x"c0",
    x"03",
    x"c0",
    x"01",
    x"80",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"01",
    x"ff",
    x"00",
    x"fe",
    x"00",
    x"fe",
    x"01",
    x"ff",
    x"f7",
    x"ff"
);
begin

process (cs)
begin
if rising_edge(cs) then
    D <= rom(to_integer(unsigned(A)));
end if;
end process;
end;

